`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 25.03.2021 17:35:43
// Design Name: 
// Module Name: GameOverPokemon
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module GameOverPokemon(
    input[6:0] X, 
    input [5:0] Y, 
    input [6:0] leftX,  
    input [5:0] topY, 
    output reg [15:0] oled_data = 16'b0
    );
    
    
    always @ (X or Y) begin
        if (X == leftX + 0 && Y == topY + 0) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 1) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 2) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 3) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 4) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 5) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 6) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 7) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 8) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 9) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 10) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 11) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 12) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 13) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 14) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 15) begin oled_data = 16'h2124; end
        else if (X == leftX + 4 && Y == topY + 15) begin oled_data = 16'h2124; end
        else if (X >= leftX + 17 && X <= leftX + 18 && Y == topY + 15) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 16) begin oled_data = 16'h2124; end
        else if (X == leftX + 4 && Y == topY + 16) begin oled_data = 16'h2124; end
        else if (X == leftX + 5 && Y == topY + 16) begin oled_data = 16'h2945; end
        else if (X == leftX + 6 && Y == topY + 16) begin oled_data = 16'h618b; end
        else if (X == leftX + 7 && Y == topY + 16) begin oled_data = 16'hbb95; end
        else if (X == leftX + 8 && Y == topY + 16) begin oled_data = 16'hbdf7; end
        else if (X == leftX + 9 && Y == topY + 16) begin oled_data = 16'hbdf7; end
        else if (X == leftX + 10 && Y == topY + 16) begin oled_data = 16'hbdf7; end
        else if (X == leftX + 11 && Y == topY + 16) begin oled_data = 16'hbdf7; end
        else if (X == leftX + 12 && Y == topY + 16) begin oled_data = 16'hbdf7; end
        else if (X == leftX + 13 && Y == topY + 16) begin oled_data = 16'hbdf7; end
        else if (X == leftX + 14 && Y == topY + 16) begin oled_data = 16'hbdf7; end
        else if (X == leftX + 15 && Y == topY + 16) begin oled_data = 16'hb5f7; end
        else if (X == leftX + 16 && Y == topY + 16) begin oled_data = 16'h3513; end
        else if (X == leftX + 17 && Y == topY + 16) begin oled_data = 16'h2a07; end
        else if (X == leftX + 37 && Y == topY + 16) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 17) begin oled_data = 16'h2124; end
        else if (X == leftX + 5 && Y == topY + 17) begin oled_data = 16'h2945; end
        else if (X == leftX + 6 && Y == topY + 17) begin oled_data = 16'h79cd; end
        else if (X == leftX + 7 && Y == topY + 17) begin oled_data = 16'hf49b; end
        else if (X == leftX + 8 && Y == topY + 17) begin oled_data = 16'hffdf; end
        else if (X >= leftX + 9 && X <= leftX + 14 && Y == topY + 17) begin oled_data = 16'hffff; end
        else if (X == leftX + 15 && Y == topY + 17) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 16 && Y == topY + 17) begin oled_data = 16'h4eda; end
        else if (X == leftX + 17 && Y == topY + 17) begin oled_data = 16'h2aca; end
        else if (X == leftX + 34 && Y == topY + 17) begin oled_data = 16'h2945; end
        else if (X == leftX + 35 && Y == topY + 17) begin oled_data = 16'h71ac; end
        else if (X == leftX + 36 && Y == topY + 17) begin oled_data = 16'hacb4; end
        else if (X == leftX + 37 && Y == topY + 17) begin oled_data = 16'had75; end
        else if (X == leftX + 38 && Y == topY + 17) begin oled_data = 16'had75; end
        else if (X == leftX + 39 && Y == topY + 17) begin oled_data = 16'ha575; end
        else if (X == leftX + 40 && Y == topY + 17) begin oled_data = 16'h33ef; end
        else if (X == leftX + 41 && Y == topY + 17) begin oled_data = 16'h2165; end
        else if (X == leftX + 0 && Y == topY + 18) begin oled_data = 16'h2124; end
        else if (X == leftX + 6 && Y == topY + 18) begin oled_data = 16'h3186; end
        else if (X == leftX + 7 && Y == topY + 18) begin oled_data = 16'h72ec; end
        else if (X == leftX + 8 && Y == topY + 18) begin oled_data = 16'hb635; end
        else if (X == leftX + 9 && Y == topY + 18) begin oled_data = 16'hbff6; end
        else if (X == leftX + 10 && Y == topY + 18) begin oled_data = 16'hbff6; end
        else if (X == leftX + 11 && Y == topY + 18) begin oled_data = 16'hbff6; end
        else if (X == leftX + 12 && Y == topY + 18) begin oled_data = 16'hbff7; end
        else if (X == leftX + 13 && Y == topY + 18) begin oled_data = 16'hef1d; end
        else if (X >= leftX + 14 && X <= leftX + 15 && Y == topY + 18) begin oled_data = 16'hffff; end
        else if (X == leftX + 16 && Y == topY + 18) begin oled_data = 16'hdfff; end
        else if (X == leftX + 17 && Y == topY + 18) begin oled_data = 16'h3638; end
        else if (X == leftX + 18 && Y == topY + 18) begin oled_data = 16'h2a27; end
        else if (X == leftX + 32 && Y == topY + 18) begin oled_data = 16'h2124; end
        else if (X == leftX + 34 && Y == topY + 18) begin oled_data = 16'h3166; end
        else if (X == leftX + 35 && Y == topY + 18) begin oled_data = 16'hb253; end
        else if (X == leftX + 36 && Y == topY + 18) begin oled_data = 16'hff3f; end
        else if (X >= leftX + 37 && X <= leftX + 39 && Y == topY + 18) begin oled_data = 16'hffff; end
        else if (X == leftX + 40 && Y == topY + 18) begin oled_data = 16'h8f7d; end
        else if (X == leftX + 41 && Y == topY + 18) begin oled_data = 16'h2a89; end
        else if (X == leftX + 48 && Y == topY + 18) begin oled_data = 16'h2945; end
        else if (X == leftX + 49 && Y == topY + 18) begin oled_data = 16'h2965; end
        else if (X == leftX + 50 && Y == topY + 18) begin oled_data = 16'h2985; end
        else if (X == leftX + 51 && Y == topY + 18) begin oled_data = 16'h29a5; end
        else if (X == leftX + 52 && Y == topY + 18) begin oled_data = 16'h2985; end
        else if (X == leftX + 57 && Y == topY + 18) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 19) begin oled_data = 16'h2124; end
        else if (X == leftX + 7 && Y == topY + 19) begin oled_data = 16'h2184; end
        else if (X == leftX + 8 && Y == topY + 19) begin oled_data = 16'h2a65; end
        else if (X == leftX + 9 && Y == topY + 19) begin oled_data = 16'h2ac5; end
        else if (X == leftX + 10 && Y == topY + 19) begin oled_data = 16'h2ac5; end
        else if (X == leftX + 11 && Y == topY + 19) begin oled_data = 16'h2ac5; end
        else if (X == leftX + 12 && Y == topY + 19) begin oled_data = 16'h630a; end
        else if (X == leftX + 13 && Y == topY + 19) begin oled_data = 16'heb9a; end
        else if (X >= leftX + 14 && X <= leftX + 15 && Y == topY + 19) begin oled_data = 16'hffff; end
        else if (X == leftX + 16 && Y == topY + 19) begin oled_data = 16'hdfff; end
        else if (X == leftX + 17 && Y == topY + 19) begin oled_data = 16'h3658; end
        else if (X == leftX + 18 && Y == topY + 19) begin oled_data = 16'h426a; end
        else if (X == leftX + 19 && Y == topY + 19) begin oled_data = 16'h9b11; end
        else if (X == leftX + 20 && Y == topY + 19) begin oled_data = 16'hb596; end
        else if (X == leftX + 21 && Y == topY + 19) begin oled_data = 16'hb596; end
        else if (X == leftX + 22 && Y == topY + 19) begin oled_data = 16'ha596; end
        else if (X == leftX + 23 && Y == topY + 19) begin oled_data = 16'h2d13; end
        else if (X == leftX + 24 && Y == topY + 19) begin oled_data = 16'h21a5; end
        else if (X == leftX + 25 && Y == topY + 19) begin oled_data = 16'h3166; end
        else if (X == leftX + 26 && Y == topY + 19) begin oled_data = 16'h822e; end
        else if (X == leftX + 27 && Y == topY + 19) begin oled_data = 16'hb596; end
        else if (X == leftX + 28 && Y == topY + 19) begin oled_data = 16'hb596; end
        else if (X == leftX + 29 && Y == topY + 19) begin oled_data = 16'hb596; end
        else if (X == leftX + 30 && Y == topY + 19) begin oled_data = 16'h4d96; end
        else if (X == leftX + 31 && Y == topY + 19) begin oled_data = 16'h2248; end
        else if (X == leftX + 34 && Y == topY + 19) begin oled_data = 16'h59aa; end
        else if (X == leftX + 35 && Y == topY + 19) begin oled_data = 16'hf47c; end
        else if (X >= leftX + 36 && X <= leftX + 37 && Y == topY + 19) begin oled_data = 16'hffff; end
        else if (X == leftX + 38 && Y == topY + 19) begin oled_data = 16'he7ff; end
        else if (X == leftX + 39 && Y == topY + 19) begin oled_data = 16'hffff; end
        else if (X == leftX + 40 && Y == topY + 19) begin oled_data = 16'hafbe; end
        else if (X == leftX + 41 && Y == topY + 19) begin oled_data = 16'h2b6c; end
        else if (X == leftX + 46 && Y == topY + 19) begin oled_data = 16'h3967; end
        else if (X == leftX + 47 && Y == topY + 19) begin oled_data = 16'hba74; end
        else if (X == leftX + 48 && Y == topY + 19) begin oled_data = 16'he67b; end
        else if (X == leftX + 49 && Y == topY + 19) begin oled_data = 16'hf77e; end
        else if (X == leftX + 50 && Y == topY + 19) begin oled_data = 16'hf7be; end
        else if (X == leftX + 51 && Y == topY + 19) begin oled_data = 16'hf7be; end
        else if (X == leftX + 52 && Y == topY + 19) begin oled_data = 16'he79e; end
        else if (X == leftX + 53 && Y == topY + 19) begin oled_data = 16'hb6fb; end
        else if (X == leftX + 54 && Y == topY + 19) begin oled_data = 16'h5d54; end
        else if (X == leftX + 55 && Y == topY + 19) begin oled_data = 16'h22aa; end
        else if (X == leftX + 0 && Y == topY + 20) begin oled_data = 16'h2124; end
        else if (X == leftX + 12 && Y == topY + 20) begin oled_data = 16'h61ab; end
        else if (X == leftX + 13 && Y == topY + 20) begin oled_data = 16'hf35a; end
        else if (X >= leftX + 14 && X <= leftX + 15 && Y == topY + 20) begin oled_data = 16'hffff; end
        else if (X == leftX + 16 && Y == topY + 20) begin oled_data = 16'hdfff; end
        else if (X == leftX + 17 && Y == topY + 20) begin oled_data = 16'h3658; end
        else if (X == leftX + 18 && Y == topY + 20) begin oled_data = 16'h428b; end
        else if (X == leftX + 19 && Y == topY + 20) begin oled_data = 16'hb394; end
        else if (X == leftX + 20 && Y == topY + 20) begin oled_data = 16'hff7e; end
        else if (X >= leftX + 21 && X <= leftX + 22 && Y == topY + 20) begin oled_data = 16'hffff; end
        else if (X == leftX + 23 && Y == topY + 20) begin oled_data = 16'h9fbe; end
        else if (X == leftX + 24 && Y == topY + 20) begin oled_data = 16'h2c91; end
        else if (X == leftX + 25 && Y == topY + 20) begin oled_data = 16'h39c8; end
        else if (X == leftX + 26 && Y == topY + 20) begin oled_data = 16'hab13; end
        else if (X == leftX + 27 && Y == topY + 20) begin oled_data = 16'hff7f; end
        else if (X >= leftX + 28 && X <= leftX + 29 && Y == topY + 20) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 20) begin oled_data = 16'hafdf; end
        else if (X == leftX + 31 && Y == topY + 20) begin oled_data = 16'h3513; end
        else if (X == leftX + 32 && Y == topY + 20) begin oled_data = 16'h2185; end
        else if (X == leftX + 34 && Y == topY + 20) begin oled_data = 16'h61aa; end
        else if (X == leftX + 35 && Y == topY + 20) begin oled_data = 16'hf4bc; end
        else if (X >= leftX + 36 && X <= leftX + 37 && Y == topY + 20) begin oled_data = 16'hffff; end
        else if (X == leftX + 38 && Y == topY + 20) begin oled_data = 16'ha73f; end
        else if (X == leftX + 39 && Y == topY + 20) begin oled_data = 16'hffdf; end
        else if (X == leftX + 40 && Y == topY + 20) begin oled_data = 16'hffff; end
        else if (X == leftX + 41 && Y == topY + 20) begin oled_data = 16'h66ba; end
        else if (X == leftX + 42 && Y == topY + 20) begin oled_data = 16'h2207; end
        else if (X == leftX + 46 && Y == topY + 20) begin oled_data = 16'h3166; end
        else if (X == leftX + 47 && Y == topY + 20) begin oled_data = 16'ha312; end
        else if (X == leftX + 48 && Y == topY + 20) begin oled_data = 16'hfdfd; end
        else if (X >= leftX + 49 && X <= leftX + 54 && Y == topY + 20) begin oled_data = 16'hffff; end
        else if (X == leftX + 55 && Y == topY + 20) begin oled_data = 16'hb7be; end
        else if (X == leftX + 56 && Y == topY + 20) begin oled_data = 16'h6d54; end
        else if (X == leftX + 57 && Y == topY + 20) begin oled_data = 16'h230b; end
        else if (X == leftX + 59 && Y == topY + 20) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 21) begin oled_data = 16'h2124; end
        else if (X == leftX + 6 && Y == topY + 21) begin oled_data = 16'h2945; end
        else if (X == leftX + 7 && Y == topY + 21) begin oled_data = 16'h618a; end
        else if (X == leftX + 8 && Y == topY + 21) begin oled_data = 16'hc355; end
        else if (X == leftX + 9 && Y == topY + 21) begin oled_data = 16'hce79; end
        else if (X == leftX + 10 && Y == topY + 21) begin oled_data = 16'hce79; end
        else if (X == leftX + 11 && Y == topY + 21) begin oled_data = 16'hce79; end
        else if (X == leftX + 12 && Y == topY + 21) begin oled_data = 16'hde9b; end
        else if (X == leftX + 13 && Y == topY + 21) begin oled_data = 16'hf6fe; end
        else if (X >= leftX + 14 && X <= leftX + 15 && Y == topY + 21) begin oled_data = 16'hffff; end
        else if (X == leftX + 16 && Y == topY + 21) begin oled_data = 16'hd7ff; end
        else if (X == leftX + 17 && Y == topY + 21) begin oled_data = 16'h3637; end
        else if (X == leftX + 18 && Y == topY + 21) begin oled_data = 16'h3228; end
        else if (X == leftX + 19 && Y == topY + 21) begin oled_data = 16'h79ed; end
        else if (X == leftX + 20 && Y == topY + 21) begin oled_data = 16'hfe7d; end
        else if (X >= leftX + 21 && X <= leftX + 23 && Y == topY + 21) begin oled_data = 16'hffff; end
        else if (X == leftX + 24 && Y == topY + 21) begin oled_data = 16'h67de; end
        else if (X == leftX + 25 && Y == topY + 21) begin oled_data = 16'h332d; end
        else if (X == leftX + 26 && Y == topY + 21) begin oled_data = 16'h9a30; end
        else if (X == leftX + 27 && Y == topY + 21) begin oled_data = 16'hff5f; end
        else if (X >= leftX + 28 && X <= leftX + 29 && Y == topY + 21) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 21) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 31 && Y == topY + 21) begin oled_data = 16'h477d; end
        else if (X == leftX + 32 && Y == topY + 21) begin oled_data = 16'h2228; end
        else if (X == leftX + 34 && Y == topY + 21) begin oled_data = 16'h69cb; end
        else if (X == leftX + 35 && Y == topY + 21) begin oled_data = 16'hfd1c; end
        else if (X >= leftX + 36 && X <= leftX + 37 && Y == topY + 21) begin oled_data = 16'hffff; end
        else if (X == leftX + 38 && Y == topY + 21) begin oled_data = 16'h8e5d; end
        else if (X == leftX + 39 && Y == topY + 21) begin oled_data = 16'hfdbd; end
        else if (X == leftX + 40 && Y == topY + 21) begin oled_data = 16'hffff; end
        else if (X == leftX + 41 && Y == topY + 21) begin oled_data = 16'hdfff; end
        else if (X == leftX + 42 && Y == topY + 21) begin oled_data = 16'h3cd2; end
        else if (X == leftX + 43 && Y == topY + 21) begin oled_data = 16'h2165; end
        else if (X == leftX + 47 && Y == topY + 21) begin oled_data = 16'h31c6; end
        else if (X == leftX + 48 && Y == topY + 21) begin oled_data = 16'h83ee; end
        else if (X == leftX + 49 && Y == topY + 21) begin oled_data = 16'h8791; end
        else if (X == leftX + 50 && Y == topY + 21) begin oled_data = 16'h5ecb; end
        else if (X == leftX + 51 && Y == topY + 21) begin oled_data = 16'h5629; end
        else if (X == leftX + 52 && Y == topY + 21) begin oled_data = 16'h85ce; end
        else if (X == leftX + 53 && Y == topY + 21) begin oled_data = 16'he55a; end
        else if (X == leftX + 54 && Y == topY + 21) begin oled_data = 16'hff7f; end
        else if (X == leftX + 55 && Y == topY + 21) begin oled_data = 16'hffff; end
        else if (X == leftX + 56 && Y == topY + 21) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 57 && Y == topY + 21) begin oled_data = 16'h677d; end
        else if (X == leftX + 58 && Y == topY + 21) begin oled_data = 16'h22ca; end
        else if (X == leftX + 60 && Y == topY + 21) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 22) begin oled_data = 16'h2124; end
        else if (X == leftX + 6 && Y == topY + 22) begin oled_data = 16'h51a9; end
        else if (X == leftX + 7 && Y == topY + 22) begin oled_data = 16'he2b9; end
        else if (X == leftX + 8 && Y == topY + 22) begin oled_data = 16'hffbf; end
        else if (X >= leftX + 9 && X <= leftX + 14 && Y == topY + 22) begin oled_data = 16'hffff; end
        else if (X == leftX + 15 && Y == topY + 22) begin oled_data = 16'hefff; end
        else if (X == leftX + 16 && Y == topY + 22) begin oled_data = 16'h475b; end
        else if (X == leftX + 17 && Y == topY + 22) begin oled_data = 16'h2b0a; end
        else if (X == leftX + 18 && Y == topY + 22) begin oled_data = 16'h2965; end
        else if (X == leftX + 19 && Y == topY + 22) begin oled_data = 16'h81ee; end
        else if (X == leftX + 20 && Y == topY + 22) begin oled_data = 16'hfebe; end
        else if (X == leftX + 21 && Y == topY + 22) begin oled_data = 16'hffff; end
        else if (X == leftX + 22 && Y == topY + 22) begin oled_data = 16'hcfff; end
        else if (X == leftX + 23 && Y == topY + 22) begin oled_data = 16'hffff; end
        else if (X == leftX + 24 && Y == topY + 22) begin oled_data = 16'ha7ff; end
        else if (X == leftX + 25 && Y == topY + 22) begin oled_data = 16'h4515; end
        else if (X == leftX + 26 && Y == topY + 22) begin oled_data = 16'hc397; end
        else if (X == leftX + 27 && Y == topY + 22) begin oled_data = 16'hffff; end
        else if (X == leftX + 28 && Y == topY + 22) begin oled_data = 16'hdfff; end
        else if (X == leftX + 29 && Y == topY + 22) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 30 && Y == topY + 22) begin oled_data = 16'hffff; end
        else if (X == leftX + 31 && Y == topY + 22) begin oled_data = 16'h4fbe; end
        else if (X == leftX + 32 && Y == topY + 22) begin oled_data = 16'h2269; end
        else if (X == leftX + 34 && Y == topY + 22) begin oled_data = 16'h51c9; end
        else if (X == leftX + 35 && Y == topY + 22) begin oled_data = 16'he439; end
        else if (X == leftX + 36 && Y == topY + 22) begin oled_data = 16'hffdf; end
        else if (X == leftX + 37 && Y == topY + 22) begin oled_data = 16'hffff; end
        else if (X == leftX + 38 && Y == topY + 22) begin oled_data = 16'h975d; end
        else if (X == leftX + 39 && Y == topY + 22) begin oled_data = 16'h9cd4; end
        else if (X == leftX + 40 && Y == topY + 22) begin oled_data = 16'hf5fc; end
        else if (X == leftX + 41 && Y == topY + 22) begin oled_data = 16'hffff; end
        else if (X == leftX + 42 && Y == topY + 22) begin oled_data = 16'hc79d; end
        else if (X == leftX + 43 && Y == topY + 22) begin oled_data = 16'h4491; end
        else if (X == leftX + 44 && Y == topY + 22) begin oled_data = 16'h2185; end
        else if (X == leftX + 48 && Y == topY + 22) begin oled_data = 16'h2184; end
        else if (X == leftX + 49 && Y == topY + 22) begin oled_data = 16'h21c4; end
        else if (X == leftX + 50 && Y == topY + 22) begin oled_data = 16'h2164; end
        else if (X == leftX + 52 && Y == topY + 22) begin oled_data = 16'h2164; end
        else if (X == leftX + 53 && Y == topY + 22) begin oled_data = 16'h5a0a; end
        else if (X == leftX + 54 && Y == topY + 22) begin oled_data = 16'heb5a; end
        else if (X == leftX + 55 && Y == topY + 22) begin oled_data = 16'hffdf; end
        else if (X == leftX + 56 && Y == topY + 22) begin oled_data = 16'hffff; end
        else if (X == leftX + 57 && Y == topY + 22) begin oled_data = 16'hc7ff; end
        else if (X == leftX + 58 && Y == topY + 22) begin oled_data = 16'h2db6; end
        else if (X == leftX + 59 && Y == topY + 22) begin oled_data = 16'h2185; end
        else if (X == leftX + 60 && Y == topY + 22) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 23) begin oled_data = 16'h2124; end
        else if (X == leftX + 6 && Y == topY + 23) begin oled_data = 16'h41a7; end
        else if (X == leftX + 7 && Y == topY + 23) begin oled_data = 16'h9bb0; end
        else if (X == leftX + 8 && Y == topY + 23) begin oled_data = 16'ha7d4; end
        else if (X == leftX + 9 && Y == topY + 23) begin oled_data = 16'ha7d4; end
        else if (X == leftX + 10 && Y == topY + 23) begin oled_data = 16'ha7d4; end
        else if (X == leftX + 11 && Y == topY + 23) begin oled_data = 16'hafd4; end
        else if (X == leftX + 12 && Y == topY + 23) begin oled_data = 16'he69b; end
        else if (X >= leftX + 13 && X <= leftX + 14 && Y == topY + 23) begin oled_data = 16'hffff; end
        else if (X == leftX + 15 && Y == topY + 23) begin oled_data = 16'hefff; end
        else if (X == leftX + 16 && Y == topY + 23) begin oled_data = 16'h3eba; end
        else if (X == leftX + 17 && Y == topY + 23) begin oled_data = 16'h2a69; end
        else if (X == leftX + 18 && Y == topY + 23) begin oled_data = 16'h3145; end
        else if (X == leftX + 19 && Y == topY + 23) begin oled_data = 16'h8a0f; end
        else if (X == leftX + 20 && Y == topY + 23) begin oled_data = 16'hff1e; end
        else if (X == leftX + 21 && Y == topY + 23) begin oled_data = 16'hffff; end
        else if (X == leftX + 22 && Y == topY + 23) begin oled_data = 16'h9fff; end
        else if (X == leftX + 23 && Y == topY + 23) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 24 && Y == topY + 23) begin oled_data = 16'hdfff; end
        else if (X == leftX + 25 && Y == topY + 23) begin oled_data = 16'h56dc; end
        else if (X == leftX + 26 && Y == topY + 23) begin oled_data = 16'he57b; end
        else if (X == leftX + 27 && Y == topY + 23) begin oled_data = 16'hffff; end
        else if (X == leftX + 28 && Y == topY + 23) begin oled_data = 16'hafff; end
        else if (X == leftX + 29 && Y == topY + 23) begin oled_data = 16'hefff; end
        else if (X == leftX + 30 && Y == topY + 23) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 31 && Y == topY + 23) begin oled_data = 16'h57be; end
        else if (X == leftX + 32 && Y == topY + 23) begin oled_data = 16'h22a9; end
        else if (X == leftX + 34 && Y == topY + 23) begin oled_data = 16'h3986; end
        else if (X == leftX + 35 && Y == topY + 23) begin oled_data = 16'hd276; end
        else if (X == leftX + 36 && Y == topY + 23) begin oled_data = 16'hffdf; end
        else if (X == leftX + 37 && Y == topY + 23) begin oled_data = 16'hffff; end
        else if (X == leftX + 38 && Y == topY + 23) begin oled_data = 16'hc7df; end
        else if (X == leftX + 39 && Y == topY + 23) begin oled_data = 16'h6c92; end
        else if (X == leftX + 40 && Y == topY + 23) begin oled_data = 16'hc396; end
        else if (X == leftX + 41 && Y == topY + 23) begin oled_data = 16'hff9f; end
        else if (X == leftX + 42 && Y == topY + 23) begin oled_data = 16'hffff; end
        else if (X == leftX + 43 && Y == topY + 23) begin oled_data = 16'hb7be; end
        else if (X == leftX + 44 && Y == topY + 23) begin oled_data = 16'h2b8d; end
        else if (X == leftX + 46 && Y == topY + 23) begin oled_data = 16'h2924; end
        else if (X == leftX + 47 && Y == topY + 23) begin oled_data = 16'h3947; end
        else if (X == leftX + 48 && Y == topY + 23) begin oled_data = 16'h4208; end
        else if (X == leftX + 49 && Y == topY + 23) begin oled_data = 16'h4228; end
        else if (X == leftX + 50 && Y == topY + 23) begin oled_data = 16'h4228; end
        else if (X == leftX + 51 && Y == topY + 23) begin oled_data = 16'h4228; end
        else if (X == leftX + 52 && Y == topY + 23) begin oled_data = 16'h2a48; end
        else if (X == leftX + 53 && Y == topY + 23) begin oled_data = 16'h3186; end
        else if (X == leftX + 54 && Y == topY + 23) begin oled_data = 16'ha992; end
        else if (X == leftX + 55 && Y == topY + 23) begin oled_data = 16'hfe5e; end
        else if (X == leftX + 56 && Y == topY + 23) begin oled_data = 16'hffff; end
        else if (X == leftX + 57 && Y == topY + 23) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 58 && Y == topY + 23) begin oled_data = 16'h471b; end
        else if (X == leftX + 59 && Y == topY + 23) begin oled_data = 16'h2207; end
        else if (X == leftX + 60 && Y == topY + 23) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 24) begin oled_data = 16'h2124; end
        else if (X == leftX + 7 && Y == topY + 24) begin oled_data = 16'h21a4; end
        else if (X == leftX + 8 && Y == topY + 24) begin oled_data = 16'h2a24; end
        else if (X == leftX + 9 && Y == topY + 24) begin oled_data = 16'h2a24; end
        else if (X == leftX + 10 && Y == topY + 24) begin oled_data = 16'h2a25; end
        else if (X == leftX + 11 && Y == topY + 24) begin oled_data = 16'h4267; end
        else if (X == leftX + 12 && Y == topY + 24) begin oled_data = 16'hab32; end
        else if (X == leftX + 13 && Y == topY + 24) begin oled_data = 16'hf63d; end
        else if (X == leftX + 14 && Y == topY + 24) begin oled_data = 16'hffff; end
        else if (X == leftX + 15 && Y == topY + 24) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 16 && Y == topY + 24) begin oled_data = 16'h8f5c; end
        else if (X == leftX + 17 && Y == topY + 24) begin oled_data = 16'h3450; end
        else if (X == leftX + 18 && Y == topY + 24) begin oled_data = 16'h622c; end
        else if (X == leftX + 19 && Y == topY + 24) begin oled_data = 16'hed7b; end
        else if (X == leftX + 20 && Y == topY + 24) begin oled_data = 16'hffff; end
        else if (X == leftX + 21 && Y == topY + 24) begin oled_data = 16'hc7ff; end
        else if (X == leftX + 22 && Y == topY + 24) begin oled_data = 16'h97bf; end
        else if (X == leftX + 23 && Y == topY + 24) begin oled_data = 16'hffff; end
        else if (X == leftX + 24 && Y == topY + 24) begin oled_data = 16'h97ff; end
        else if (X == leftX + 25 && Y == topY + 24) begin oled_data = 16'haf3e; end
        else if (X == leftX + 26 && Y == topY + 24) begin oled_data = 16'hffdf; end
        else if (X == leftX + 27 && Y == topY + 24) begin oled_data = 16'hb7ff; end
        else if (X == leftX + 28 && Y == topY + 24) begin oled_data = 16'hafff; end
        else if (X == leftX + 29 && Y == topY + 24) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 24) begin oled_data = 16'hafff; end
        else if (X == leftX + 31 && Y == topY + 24) begin oled_data = 16'h3594; end
        else if (X == leftX + 32 && Y == topY + 24) begin oled_data = 16'h2165; end
        else if (X == leftX + 33 && Y == topY + 24) begin oled_data = 16'h2944; end
        else if (X == leftX + 34 && Y == topY + 24) begin oled_data = 16'h69ac; end
        else if (X == leftX + 35 && Y == topY + 24) begin oled_data = 16'hecdb; end
        else if (X >= leftX + 36 && X <= leftX + 42 && Y == topY + 24) begin oled_data = 16'hffff; end
        else if (X == leftX + 43 && Y == topY + 24) begin oled_data = 16'he7ff; end
        else if (X == leftX + 44 && Y == topY + 24) begin oled_data = 16'h3d13; end
        else if (X == leftX + 45 && Y == topY + 24) begin oled_data = 16'h2985; end
        else if (X == leftX + 46 && Y == topY + 24) begin oled_data = 16'h916f; end
        else if (X == leftX + 47 && Y == topY + 24) begin oled_data = 16'hf53c; end
        else if (X == leftX + 48 && Y == topY + 24) begin oled_data = 16'hffdf; end
        else if (X >= leftX + 49 && X <= leftX + 50 && Y == topY + 24) begin oled_data = 16'hffff; end
        else if (X == leftX + 51 && Y == topY + 24) begin oled_data = 16'hb7ff; end
        else if (X == leftX + 52 && Y == topY + 24) begin oled_data = 16'h3e16; end
        else if (X == leftX + 53 && Y == topY + 24) begin oled_data = 16'h5a0c; end
        else if (X == leftX + 54 && Y == topY + 24) begin oled_data = 16'heb5a; end
        else if (X == leftX + 55 && Y == topY + 24) begin oled_data = 16'hff9f; end
        else if (X == leftX + 56 && Y == topY + 24) begin oled_data = 16'hffff; end
        else if (X == leftX + 57 && Y == topY + 24) begin oled_data = 16'h9fff; end
        else if (X == leftX + 58 && Y == topY + 24) begin oled_data = 16'h3512; end
        else if (X == leftX + 59 && Y == topY + 24) begin oled_data = 16'h2185; end
        else if (X == leftX + 60 && Y == topY + 24) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 25) begin oled_data = 16'h2124; end
        else if (X == leftX + 11 && Y == topY + 25) begin oled_data = 16'h3146; end
        else if (X == leftX + 12 && Y == topY + 25) begin oled_data = 16'h89ee; end
        else if (X == leftX + 13 && Y == topY + 25) begin oled_data = 16'hec9b; end
        else if (X >= leftX + 14 && X <= leftX + 15 && Y == topY + 25) begin oled_data = 16'hffff; end
        else if (X == leftX + 16 && Y == topY + 25) begin oled_data = 16'hb7df; end
        else if (X == leftX + 17 && Y == topY + 25) begin oled_data = 16'h3db5; end
        else if (X == leftX + 18 && Y == topY + 25) begin oled_data = 16'h6a8e; end
        else if (X == leftX + 19 && Y == topY + 25) begin oled_data = 16'hf5fd; end
        else if (X == leftX + 20 && Y == topY + 25) begin oled_data = 16'hffff; end
        else if (X == leftX + 21 && Y == topY + 25) begin oled_data = 16'hbfff; end
        else if (X == leftX + 22 && Y == topY + 25) begin oled_data = 16'h865d; end
        else if (X == leftX + 23 && Y == topY + 25) begin oled_data = 16'hffdf; end
        else if (X == leftX + 24 && Y == topY + 25) begin oled_data = 16'hc7ff; end
        else if (X == leftX + 25 && Y == topY + 25) begin oled_data = 16'hc7ff; end
        else if (X == leftX + 26 && Y == topY + 25) begin oled_data = 16'hffff; end
        else if (X == leftX + 27 && Y == topY + 25) begin oled_data = 16'h7fdf; end
        else if (X == leftX + 28 && Y == topY + 25) begin oled_data = 16'hcefe; end
        else if (X == leftX + 29 && Y == topY + 25) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 25) begin oled_data = 16'hb7ff; end
        else if (X == leftX + 31 && Y == topY + 25) begin oled_data = 16'h2d54; end
        else if (X == leftX + 32 && Y == topY + 25) begin oled_data = 16'h2165; end
        else if (X == leftX + 33 && Y == topY + 25) begin oled_data = 16'h4187; end
        else if (X == leftX + 34 && Y == topY + 25) begin oled_data = 16'hcb16; end
        else if (X == leftX + 35 && Y == topY + 25) begin oled_data = 16'hffdf; end
        else if (X == leftX + 36 && Y == topY + 25) begin oled_data = 16'hffff; end
        else if (X == leftX + 37 && Y == topY + 25) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 38 && Y == topY + 25) begin oled_data = 16'hc7fb; end
        else if (X == leftX + 39 && Y == topY + 25) begin oled_data = 16'hc7d7; end
        else if (X == leftX + 40 && Y == topY + 25) begin oled_data = 16'hcf99; end
        else if (X == leftX + 41 && Y == topY + 25) begin oled_data = 16'hff5e; end
        else if (X == leftX + 42 && Y == topY + 25) begin oled_data = 16'hffff; end
        else if (X == leftX + 43 && Y == topY + 25) begin oled_data = 16'hdfff; end
        else if (X == leftX + 44 && Y == topY + 25) begin oled_data = 16'h4d33; end
        else if (X == leftX + 45 && Y == topY + 25) begin oled_data = 16'h29a6; end
        else if (X == leftX + 46 && Y == topY + 25) begin oled_data = 16'ha191; end
        else if (X == leftX + 47 && Y == topY + 25) begin oled_data = 16'hfdde; end
        else if (X >= leftX + 48 && X <= leftX + 49 && Y == topY + 25) begin oled_data = 16'hffff; end
        else if (X == leftX + 50 && Y == topY + 25) begin oled_data = 16'hdffc; end
        else if (X == leftX + 51 && Y == topY + 25) begin oled_data = 16'h97fb; end
        else if (X == leftX + 52 && Y == topY + 25) begin oled_data = 16'h34d1; end
        else if (X == leftX + 53 && Y == topY + 25) begin oled_data = 16'h69ac; end
        else if (X == leftX + 54 && Y == topY + 25) begin oled_data = 16'hfc1c; end
        else if (X >= leftX + 55 && X <= leftX + 56 && Y == topY + 25) begin oled_data = 16'hffff; end
        else if (X == leftX + 57 && Y == topY + 25) begin oled_data = 16'h7fff; end
        else if (X == leftX + 58 && Y == topY + 25) begin oled_data = 16'h2bad; end
        else if (X == leftX + 0 && Y == topY + 26) begin oled_data = 16'h2124; end
        else if (X == leftX + 4 && Y == topY + 26) begin oled_data = 16'h2124; end
        else if (X == leftX + 5 && Y == topY + 26) begin oled_data = 16'h2944; end
        else if (X == leftX + 6 && Y == topY + 26) begin oled_data = 16'h5188; end
        else if (X == leftX + 7 && Y == topY + 26) begin oled_data = 16'h8acf; end
        else if (X == leftX + 8 && Y == topY + 26) begin oled_data = 16'h9492; end
        else if (X == leftX + 9 && Y == topY + 26) begin oled_data = 16'h94b2; end
        else if (X == leftX + 10 && Y == topY + 26) begin oled_data = 16'h94b2; end
        else if (X == leftX + 11 && Y == topY + 26) begin oled_data = 16'hacf4; end
        else if (X == leftX + 12 && Y == topY + 26) begin oled_data = 16'hf59c; end
        else if (X >= leftX + 13 && X <= leftX + 14 && Y == topY + 26) begin oled_data = 16'hffff; end
        else if (X == leftX + 15 && Y == topY + 26) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 16 && Y == topY + 26) begin oled_data = 16'h6f7c; end
        else if (X == leftX + 17 && Y == topY + 26) begin oled_data = 16'h344f; end
        else if (X == leftX + 18 && Y == topY + 26) begin oled_data = 16'h41e8; end
        else if (X == leftX + 19 && Y == topY + 26) begin oled_data = 16'hbbb4; end
        else if (X == leftX + 20 && Y == topY + 26) begin oled_data = 16'hffdf; end
        else if (X == leftX + 21 && Y == topY + 26) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 22 && Y == topY + 26) begin oled_data = 16'h779f; end
        else if (X == leftX + 23 && Y == topY + 26) begin oled_data = 16'hae38; end
        else if (X == leftX + 24 && Y == topY + 26) begin oled_data = 16'hf7df; end
        else if (X == leftX + 25 && Y == topY + 26) begin oled_data = 16'hefff; end
        else if (X == leftX + 26 && Y == topY + 26) begin oled_data = 16'hffff; end
        else if (X == leftX + 27 && Y == topY + 26) begin oled_data = 16'hb7ff; end
        else if (X == leftX + 28 && Y == topY + 26) begin oled_data = 16'h865c; end
        else if (X == leftX + 29 && Y == topY + 26) begin oled_data = 16'hff5e; end
        else if (X == leftX + 30 && Y == topY + 26) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 31 && Y == topY + 26) begin oled_data = 16'h777d; end
        else if (X == leftX + 32 && Y == topY + 26) begin oled_data = 16'h2b6d; end
        else if (X == leftX + 33 && Y == topY + 26) begin oled_data = 16'h5189; end
        else if (X == leftX + 34 && Y == topY + 26) begin oled_data = 16'hcbb7; end
        else if (X == leftX + 35 && Y == topY + 26) begin oled_data = 16'hffbf; end
        else if (X == leftX + 36 && Y == topY + 26) begin oled_data = 16'hffff; end
        else if (X == leftX + 37 && Y == topY + 26) begin oled_data = 16'hc7be; end
        else if (X == leftX + 38 && Y == topY + 26) begin oled_data = 16'h3cb1; end
        else if (X == leftX + 39 && Y == topY + 26) begin oled_data = 16'h2a05; end
        else if (X == leftX + 40 && Y == topY + 26) begin oled_data = 16'h4a68; end
        else if (X == leftX + 41 && Y == topY + 26) begin oled_data = 16'hdbb8; end
        else if (X >= leftX + 42 && X <= leftX + 43 && Y == topY + 26) begin oled_data = 16'hffff; end
        else if (X == leftX + 44 && Y == topY + 26) begin oled_data = 16'ha7be; end
        else if (X == leftX + 45 && Y == topY + 26) begin oled_data = 16'h332c; end
        else if (X == leftX + 46 && Y == topY + 26) begin oled_data = 16'h69cb; end
        else if (X == leftX + 47 && Y == topY + 26) begin oled_data = 16'hec3a; end
        else if (X == leftX + 48 && Y == topY + 26) begin oled_data = 16'hffbf; end
        else if (X == leftX + 49 && Y == topY + 26) begin oled_data = 16'hefff; end
        else if (X == leftX + 50 && Y == topY + 26) begin oled_data = 16'h77d7; end
        else if (X == leftX + 51 && Y == topY + 26) begin oled_data = 16'h360d; end
        else if (X == leftX + 52 && Y == topY + 26) begin oled_data = 16'h29e5; end
        else if (X == leftX + 53 && Y == topY + 26) begin oled_data = 16'h618b; end
        else if (X == leftX + 54 && Y == topY + 26) begin oled_data = 16'hebda; end
        else if (X == leftX + 55 && Y == topY + 26) begin oled_data = 16'hffdf; end
        else if (X == leftX + 56 && Y == topY + 26) begin oled_data = 16'hffff; end
        else if (X == leftX + 57 && Y == topY + 26) begin oled_data = 16'hafff; end
        else if (X == leftX + 58 && Y == topY + 26) begin oled_data = 16'h2d13; end
        else if (X == leftX + 59 && Y == topY + 26) begin oled_data = 16'h2185; end
        else if (X == leftX + 0 && Y == topY + 27) begin oled_data = 16'h2124; end
        else if (X == leftX + 6 && Y == topY + 27) begin oled_data = 16'h4988; end
        else if (X == leftX + 7 && Y == topY + 27) begin oled_data = 16'hc295; end
        else if (X == leftX + 8 && Y == topY + 27) begin oled_data = 16'hff3f; end
        else if (X >= leftX + 9 && X <= leftX + 15 && Y == topY + 27) begin oled_data = 16'hffff; end
        else if (X == leftX + 16 && Y == topY + 27) begin oled_data = 16'hcfff; end
        else if (X == leftX + 17 && Y == topY + 27) begin oled_data = 16'h3e38; end
        else if (X == leftX + 18 && Y == topY + 27) begin oled_data = 16'h6a8e; end
        else if (X == leftX + 19 && Y == topY + 27) begin oled_data = 16'he59b; end
        else if (X == leftX + 20 && Y == topY + 27) begin oled_data = 16'hffff; end
        else if (X == leftX + 21 && Y == topY + 27) begin oled_data = 16'hc7ff; end
        else if (X == leftX + 22 && Y == topY + 27) begin oled_data = 16'h56da; end
        else if (X == leftX + 23 && Y == topY + 27) begin oled_data = 16'hccd9; end
        else if (X == leftX + 24 && Y == topY + 27) begin oled_data = 16'hffdf; end
        else if (X == leftX + 25 && Y == topY + 27) begin oled_data = 16'hffff; end
        else if (X == leftX + 26 && Y == topY + 27) begin oled_data = 16'hdfff; end
        else if (X == leftX + 27 && Y == topY + 27) begin oled_data = 16'h5f7c; end
        else if (X == leftX + 28 && Y == topY + 27) begin oled_data = 16'hc57a; end
        else if (X == leftX + 29 && Y == topY + 27) begin oled_data = 16'hffbf; end
        else if (X == leftX + 30 && Y == topY + 27) begin oled_data = 16'hdfff; end
        else if (X == leftX + 31 && Y == topY + 27) begin oled_data = 16'h471a; end
        else if (X == leftX + 32 && Y == topY + 27) begin oled_data = 16'h3289; end
        else if (X == leftX + 33 && Y == topY + 27) begin oled_data = 16'h9a30; end
        else if (X == leftX + 34 && Y == topY + 27) begin oled_data = 16'hfe9e; end
        else if (X >= leftX + 35 && X <= leftX + 36 && Y == topY + 27) begin oled_data = 16'hffff; end
        else if (X == leftX + 37 && Y == topY + 27) begin oled_data = 16'h5e99; end
        else if (X == leftX + 38 && Y == topY + 27) begin oled_data = 16'h29e7; end
        else if (X == leftX + 40 && Y == topY + 27) begin oled_data = 16'h49c8; end
        else if (X == leftX + 41 && Y == topY + 27) begin oled_data = 16'hd437; end
        else if (X == leftX + 42 && Y == topY + 27) begin oled_data = 16'hff9f; end
        else if (X == leftX + 43 && Y == topY + 27) begin oled_data = 16'hffff; end
        else if (X == leftX + 44 && Y == topY + 27) begin oled_data = 16'hb7be; end
        else if (X == leftX + 45 && Y == topY + 27) begin oled_data = 16'h338d; end
        else if (X == leftX + 46 && Y == topY + 27) begin oled_data = 16'h698b; end
        else if (X == leftX + 47 && Y == topY + 27) begin oled_data = 16'hdbb9; end
        else if (X == leftX + 48 && Y == topY + 27) begin oled_data = 16'hffbf; end
        else if (X == leftX + 49 && Y == topY + 27) begin oled_data = 16'hefff; end
        else if (X == leftX + 50 && Y == topY + 27) begin oled_data = 16'h77bd; end
        else if (X == leftX + 51 && Y == topY + 27) begin oled_data = 16'h3bcf; end
        else if (X == leftX + 52 && Y == topY + 27) begin oled_data = 16'h69ab; end
        else if (X == leftX + 53 && Y == topY + 27) begin oled_data = 16'hb3d4; end
        else if (X == leftX + 54 && Y == topY + 27) begin oled_data = 16'hf63d; end
        else if (X == leftX + 55 && Y == topY + 27) begin oled_data = 16'hffff; end
        else if (X == leftX + 56 && Y == topY + 27) begin oled_data = 16'he7ff; end
        else if (X == leftX + 57 && Y == topY + 27) begin oled_data = 16'h87d8; end
        else if (X == leftX + 58 && Y == topY + 27) begin oled_data = 16'h344f; end
        else if (X == leftX + 59 && Y == topY + 27) begin oled_data = 16'h2165; end
        else if (X == leftX + 0 && Y == topY + 28) begin oled_data = 16'h2124; end
        else if (X == leftX + 5 && Y == topY + 28) begin oled_data = 16'h3166; end
        else if (X == leftX + 6 && Y == topY + 28) begin oled_data = 16'h8a0f; end
        else if (X == leftX + 7 && Y == topY + 28) begin oled_data = 16'hd679; end
        else if (X == leftX + 8 && Y == topY + 28) begin oled_data = 16'hd7fa; end
        else if (X == leftX + 9 && Y == topY + 28) begin oled_data = 16'hd7fa; end
        else if (X == leftX + 10 && Y == topY + 28) begin oled_data = 16'hd7fa; end
        else if (X == leftX + 11 && Y == topY + 28) begin oled_data = 16'hd7fa; end
        else if (X == leftX + 12 && Y == topY + 28) begin oled_data = 16'hd7fa; end
        else if (X == leftX + 13 && Y == topY + 28) begin oled_data = 16'hd7fa; end
        else if (X == leftX + 14 && Y == topY + 28) begin oled_data = 16'hd7fa; end
        else if (X == leftX + 15 && Y == topY + 28) begin oled_data = 16'hcffa; end
        else if (X == leftX + 16 && Y == topY + 28) begin oled_data = 16'h4697; end
        else if (X == leftX + 17 && Y == topY + 28) begin oled_data = 16'h2ac9; end
        else if (X == leftX + 18 && Y == topY + 28) begin oled_data = 16'h41c8; end
        else if (X == leftX + 19 && Y == topY + 28) begin oled_data = 16'hc3d5; end
        else if (X == leftX + 20 && Y == topY + 28) begin oled_data = 16'hffff; end
        else if (X == leftX + 21 && Y == topY + 28) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 22 && Y == topY + 28) begin oled_data = 16'h5fbe; end
        else if (X == leftX + 23 && Y == topY + 28) begin oled_data = 16'h6431; end
        else if (X == leftX + 24 && Y == topY + 28) begin oled_data = 16'hd5f9; end
        else if (X == leftX + 25 && Y == topY + 28) begin oled_data = 16'hffff; end
        else if (X == leftX + 26 && Y == topY + 28) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 27 && Y == topY + 28) begin oled_data = 16'h5f9e; end
        else if (X == leftX + 28 && Y == topY + 28) begin oled_data = 16'h8413; end
        else if (X == leftX + 29 && Y == topY + 28) begin oled_data = 16'hf6dd; end
        else if (X == leftX + 30 && Y == topY + 28) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 31 && Y == topY + 28) begin oled_data = 16'h475d; end
        else if (X == leftX + 32 && Y == topY + 28) begin oled_data = 16'h2a28; end
        else if (X == leftX + 33 && Y == topY + 28) begin oled_data = 16'h5a8a; end
        else if (X == leftX + 34 && Y == topY + 28) begin oled_data = 16'ha5f2; end
        else if (X == leftX + 35 && Y == topY + 28) begin oled_data = 16'ha714; end
        else if (X == leftX + 36 && Y == topY + 28) begin oled_data = 16'ha6f4; end
        else if (X == leftX + 37 && Y == topY + 28) begin oled_data = 16'h5cd2; end
        else if (X == leftX + 38 && Y == topY + 28) begin oled_data = 16'h29c6; end
        else if (X == leftX + 40 && Y == topY + 28) begin oled_data = 16'h2164; end
        else if (X == leftX + 41 && Y == topY + 28) begin oled_data = 16'h52a9; end
        else if (X == leftX + 42 && Y == topY + 28) begin oled_data = 16'ha5b2; end
        else if (X == leftX + 43 && Y == topY + 28) begin oled_data = 16'ha714; end
        else if (X == leftX + 44 && Y == topY + 28) begin oled_data = 16'ha6f4; end
        else if (X == leftX + 45 && Y == topY + 28) begin oled_data = 16'h54b1; end
        else if (X == leftX + 46 && Y == topY + 28) begin oled_data = 16'h6a0c; end
        else if (X == leftX + 47 && Y == topY + 28) begin oled_data = 16'he3fa; end
        else if (X == leftX + 48 && Y == topY + 28) begin oled_data = 16'hffbf; end
        else if (X == leftX + 49 && Y == topY + 28) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 50 && Y == topY + 28) begin oled_data = 16'hc7bd; end
        else if (X == leftX + 51 && Y == topY + 28) begin oled_data = 16'hd65a; end
        else if (X == leftX + 52 && Y == topY + 28) begin oled_data = 16'hff3e; end
        else if (X >= leftX + 53 && X <= leftX + 55 && Y == topY + 28) begin oled_data = 16'hffff; end
        else if (X == leftX + 56 && Y == topY + 28) begin oled_data = 16'hafff; end
        else if (X == leftX + 57 && Y == topY + 28) begin oled_data = 16'h35f3; end
        else if (X == leftX + 58 && Y == topY + 28) begin oled_data = 16'h21a5; end
        else if (X == leftX + 0 && Y == topY + 29) begin oled_data = 16'h2124; end
        else if (X == leftX + 6 && Y == topY + 29) begin oled_data = 16'h29c5; end
        else if (X == leftX + 7 && Y == topY + 29) begin oled_data = 16'h3386; end
        else if (X == leftX + 8 && Y == topY + 29) begin oled_data = 16'h33c5; end
        else if (X == leftX + 9 && Y == topY + 29) begin oled_data = 16'h33c5; end
        else if (X == leftX + 10 && Y == topY + 29) begin oled_data = 16'h33c5; end
        else if (X == leftX + 11 && Y == topY + 29) begin oled_data = 16'h33c5; end
        else if (X == leftX + 12 && Y == topY + 29) begin oled_data = 16'h33c5; end
        else if (X == leftX + 13 && Y == topY + 29) begin oled_data = 16'h33c5; end
        else if (X == leftX + 14 && Y == topY + 29) begin oled_data = 16'h33c5; end
        else if (X == leftX + 15 && Y == topY + 29) begin oled_data = 16'h33a6; end
        else if (X == leftX + 16 && Y == topY + 29) begin oled_data = 16'h2a25; end
        else if (X == leftX + 17 && Y == topY + 29) begin oled_data = 16'h2965; end
        else if (X == leftX + 18 && Y == topY + 29) begin oled_data = 16'h81ed; end
        else if (X == leftX + 19 && Y == topY + 29) begin oled_data = 16'heebc; end
        else if (X == leftX + 20 && Y == topY + 29) begin oled_data = 16'hf7fe; end
        else if (X == leftX + 21 && Y == topY + 29) begin oled_data = 16'ha7fd; end
        else if (X == leftX + 22 && Y == topY + 29) begin oled_data = 16'h3d94; end
        else if (X == leftX + 23 && Y == topY + 29) begin oled_data = 16'h726d; end
        else if (X == leftX + 24 && Y == topY + 29) begin oled_data = 16'hd6b9; end
        else if (X == leftX + 25 && Y == topY + 29) begin oled_data = 16'hd7fa; end
        else if (X == leftX + 26 && Y == topY + 29) begin oled_data = 16'h779a; end
        else if (X == leftX + 27 && Y == topY + 29) begin oled_data = 16'h5490; end
        else if (X == leftX + 28 && Y == topY + 29) begin oled_data = 16'hc437; end
        else if (X == leftX + 29 && Y == topY + 29) begin oled_data = 16'hf7be; end
        else if (X == leftX + 30 && Y == topY + 29) begin oled_data = 16'hdffe; end
        else if (X == leftX + 31 && Y == topY + 29) begin oled_data = 16'h36b9; end
        else if (X == leftX + 32 && Y == topY + 29) begin oled_data = 16'h21c6; end
        else if (X == leftX + 34 && Y == topY + 29) begin oled_data = 16'h2164; end
        else if (X == leftX + 35 && Y == topY + 29) begin oled_data = 16'h2164; end
        else if (X == leftX + 36 && Y == topY + 29) begin oled_data = 16'h2164; end
        else if (X == leftX + 38 && Y == topY + 29) begin oled_data = 16'h2124; end
        else if (X == leftX + 42 && Y == topY + 29) begin oled_data = 16'h2164; end
        else if (X == leftX + 43 && Y == topY + 29) begin oled_data = 16'h2164; end
        else if (X == leftX + 44 && Y == topY + 29) begin oled_data = 16'h2164; end
        else if (X == leftX + 46 && Y == topY + 29) begin oled_data = 16'h5189; end
        else if (X == leftX + 47 && Y == topY + 29) begin oled_data = 16'hd377; end
        else if (X == leftX + 48 && Y == topY + 29) begin oled_data = 16'hff9f; end
        else if (X >= leftX + 49 && X <= leftX + 53 && Y == topY + 29) begin oled_data = 16'hffff; end
        else if (X == leftX + 54 && Y == topY + 29) begin oled_data = 16'hcffb; end
        else if (X == leftX + 55 && Y == topY + 29) begin oled_data = 16'h9ff4; end
        else if (X == leftX + 56 && Y == topY + 29) begin oled_data = 16'h46b2; end
        else if (X == leftX + 57 && Y == topY + 29) begin oled_data = 16'h2a67; end
        else if (X == leftX + 0 && Y == topY + 30) begin oled_data = 16'h2124; end
        else if (X == leftX + 18 && Y == topY + 30) begin oled_data = 16'h31c5; end
        else if (X == leftX + 19 && Y == topY + 30) begin oled_data = 16'h3be7; end
        else if (X == leftX + 20 && Y == topY + 30) begin oled_data = 16'h3c67; end
        else if (X == leftX + 21 && Y == topY + 30) begin oled_data = 16'h3407; end
        else if (X == leftX + 22 && Y == topY + 30) begin oled_data = 16'h21c5; end
        else if (X == leftX + 23 && Y == topY + 30) begin oled_data = 16'h29a5; end
        else if (X == leftX + 24 && Y == topY + 30) begin oled_data = 16'h3305; end
        else if (X == leftX + 25 && Y == topY + 30) begin oled_data = 16'h3365; end
        else if (X == leftX + 26 && Y == topY + 30) begin oled_data = 16'h2aa5; end
        else if (X == leftX + 27 && Y == topY + 30) begin oled_data = 16'h2965; end
        else if (X == leftX + 28 && Y == topY + 30) begin oled_data = 16'h3ac6; end
        else if (X == leftX + 29 && Y == topY + 30) begin oled_data = 16'h4467; end
        else if (X == leftX + 30 && Y == topY + 30) begin oled_data = 16'h3c67; end
        else if (X == leftX + 31 && Y == topY + 30) begin oled_data = 16'h2aa6; end
        else if (X == leftX + 46 && Y == topY + 30) begin oled_data = 16'h2984; end
        else if (X == leftX + 47 && Y == topY + 30) begin oled_data = 16'h4407; end
        else if (X == leftX + 48 && Y == topY + 30) begin oled_data = 16'h65eb; end
        else if (X == leftX + 49 && Y == topY + 30) begin oled_data = 16'h870e; end
        else if (X == leftX + 50 && Y == topY + 30) begin oled_data = 16'h8f90; end
        else if (X == leftX + 51 && Y == topY + 30) begin oled_data = 16'h8f90; end
        else if (X == leftX + 52 && Y == topY + 30) begin oled_data = 16'h7f6f; end
        else if (X == leftX + 53 && Y == topY + 30) begin oled_data = 16'h56cb; end
        else if (X == leftX + 54 && Y == topY + 30) begin oled_data = 16'h34e6; end
        else if (X == leftX + 55 && Y == topY + 30) begin oled_data = 16'h2ac5; end
        else if (X == leftX + 56 && Y == topY + 30) begin oled_data = 16'h21a4; end
        else if (X == leftX + 0 && Y == topY + 31) begin oled_data = 16'h2124; end
        else if (X == leftX + 26 && Y == topY + 31) begin oled_data = 16'h2124; end
        else if (X == leftX + 49 && Y == topY + 31) begin oled_data = 16'h2164; end
        else if (X == leftX + 50 && Y == topY + 31) begin oled_data = 16'h2184; end
        else if (X == leftX + 51 && Y == topY + 31) begin oled_data = 16'h2184; end
        else if (X == leftX + 52 && Y == topY + 31) begin oled_data = 16'h2184; end
        else if (X == leftX + 0 && Y == topY + 32) begin oled_data = 16'h2124; end
        else if (X == leftX + 11 && Y == topY + 32) begin oled_data = 16'h2124; end
        else if (X == leftX + 20 && Y == topY + 32) begin oled_data = 16'h2945; end
        else if (X == leftX + 21 && Y == topY + 32) begin oled_data = 16'h596a; end
        else if (X == leftX + 22 && Y == topY + 32) begin oled_data = 16'h8b70; end
        else if (X == leftX + 23 && Y == topY + 32) begin oled_data = 16'h8450; end
        else if (X == leftX + 24 && Y == topY + 32) begin oled_data = 16'h8450; end
        else if (X == leftX + 25 && Y == topY + 32) begin oled_data = 16'h8450; end
        else if (X == leftX + 26 && Y == topY + 32) begin oled_data = 16'h8450; end
        else if (X == leftX + 27 && Y == topY + 32) begin oled_data = 16'h8450; end
        else if (X == leftX + 28 && Y == topY + 32) begin oled_data = 16'h8450; end
        else if (X == leftX + 29 && Y == topY + 32) begin oled_data = 16'h8450; end
        else if (X == leftX + 30 && Y == topY + 32) begin oled_data = 16'h33ef; end
        else if (X == leftX + 31 && Y == topY + 32) begin oled_data = 16'h29c6; end
        else if (X == leftX + 38 && Y == topY + 32) begin oled_data = 16'h2124; end
        else if (X == leftX + 41 && Y == topY + 32) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 33) begin oled_data = 16'h2124; end
        else if (X >= leftX + 9 && X <= leftX + 10 && Y == topY + 33) begin oled_data = 16'h2124; end
        else if (X == leftX + 11 && Y == topY + 33) begin oled_data = 16'h3145; end
        else if (X == leftX + 12 && Y == topY + 33) begin oled_data = 16'h39c7; end
        else if (X == leftX + 13 && Y == topY + 33) begin oled_data = 16'h4248; end
        else if (X == leftX + 14 && Y == topY + 33) begin oled_data = 16'h4a69; end
        else if (X == leftX + 15 && Y == topY + 33) begin oled_data = 16'h4a89; end
        else if (X == leftX + 16 && Y == topY + 33) begin oled_data = 16'h4269; end
        else if (X == leftX + 17 && Y == topY + 33) begin oled_data = 16'h3a28; end
        else if (X == leftX + 18 && Y == topY + 33) begin oled_data = 16'h29e6; end
        else if (X == leftX + 19 && Y == topY + 33) begin oled_data = 16'h2185; end
        else if (X == leftX + 20 && Y == topY + 33) begin oled_data = 16'h3166; end
        else if (X == leftX + 21 && Y == topY + 33) begin oled_data = 16'h99d1; end
        else if (X == leftX + 22 && Y == topY + 33) begin oled_data = 16'hfe3e; end
        else if (X >= leftX + 23 && X <= leftX + 29 && Y == topY + 33) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 33) begin oled_data = 16'h573c; end
        else if (X == leftX + 31 && Y == topY + 33) begin oled_data = 16'h3aab; end
        else if (X == leftX + 32 && Y == topY + 33) begin oled_data = 16'h9a31; end
        else if (X == leftX + 33 && Y == topY + 33) begin oled_data = 16'hb3d4; end
        else if (X == leftX + 34 && Y == topY + 33) begin oled_data = 16'habd3; end
        else if (X == leftX + 35 && Y == topY + 33) begin oled_data = 16'h63cf; end
        else if (X == leftX + 36 && Y == topY + 33) begin oled_data = 16'h2a68; end
        else if (X == leftX + 37 && Y == topY + 33) begin oled_data = 16'h2165; end
        else if (X == leftX + 38 && Y == topY + 33) begin oled_data = 16'h2944; end
        else if (X == leftX + 39 && Y == topY + 33) begin oled_data = 16'h5189; end
        else if (X == leftX + 40 && Y == topY + 33) begin oled_data = 16'haa52; end
        else if (X == leftX + 41 && Y == topY + 33) begin oled_data = 16'hb3d4; end
        else if (X == leftX + 42 && Y == topY + 33) begin oled_data = 16'habd3; end
        else if (X == leftX + 43 && Y == topY + 33) begin oled_data = 16'h63af; end
        else if (X == leftX + 44 && Y == topY + 33) begin oled_data = 16'h2a07; end
        else if (X == leftX + 48 && Y == topY + 33) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 34) begin oled_data = 16'h2124; end
        else if (X == leftX + 8 && Y == topY + 34) begin oled_data = 16'h2944; end
        else if (X == leftX + 9 && Y == topY + 34) begin oled_data = 16'h5989; end
        else if (X == leftX + 10 && Y == topY + 34) begin oled_data = 16'hb374; end
        else if (X == leftX + 11 && Y == topY + 34) begin oled_data = 16'he69c; end
        else if (X == leftX + 12 && Y == topY + 34) begin oled_data = 16'hffbf; end
        else if (X >= leftX + 13 && X <= leftX + 17 && Y == topY + 34) begin oled_data = 16'hffff; end
        else if (X == leftX + 18 && Y == topY + 34) begin oled_data = 16'hb7dc; end
        else if (X == leftX + 19 && Y == topY + 34) begin oled_data = 16'h2e77; end
        else if (X == leftX + 20 && Y == topY + 34) begin oled_data = 16'h29c6; end
        else if (X == leftX + 21 && Y == topY + 34) begin oled_data = 16'h49c8; end
        else if (X == leftX + 22 && Y == topY + 34) begin oled_data = 16'habd2; end
        else if (X == leftX + 23 && Y == topY + 34) begin oled_data = 16'hdf7a; end
        else if (X == leftX + 24 && Y == topY + 34) begin oled_data = 16'hdffa; end
        else if (X == leftX + 25 && Y == topY + 34) begin oled_data = 16'hdffa; end
        else if (X == leftX + 26 && Y == topY + 34) begin oled_data = 16'hdffa; end
        else if (X == leftX + 27 && Y == topY + 34) begin oled_data = 16'hef9c; end
        else if (X == leftX + 28 && Y == topY + 34) begin oled_data = 16'hffdf; end
        else if (X == leftX + 29 && Y == topY + 34) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 34) begin oled_data = 16'hd7df; end
        else if (X == leftX + 31 && Y == topY + 34) begin oled_data = 16'h45d7; end
        else if (X == leftX + 32 && Y == topY + 34) begin oled_data = 16'h9b12; end
        else if (X == leftX + 33 && Y == topY + 34) begin oled_data = 16'hffbf; end
        else if (X == leftX + 34 && Y == topY + 34) begin oled_data = 16'hffff; end
        else if (X == leftX + 35 && Y == topY + 34) begin oled_data = 16'hd7ff; end
        else if (X == leftX + 36 && Y == topY + 34) begin oled_data = 16'h3d75; end
        else if (X == leftX + 37 && Y == topY + 34) begin oled_data = 16'h2207; end
        else if (X == leftX + 38 && Y == topY + 34) begin oled_data = 16'h2945; end
        else if (X == leftX + 39 && Y == topY + 34) begin oled_data = 16'h79cd; end
        else if (X == leftX + 40 && Y == topY + 34) begin oled_data = 16'hed5c; end
        else if (X >= leftX + 41 && X <= leftX + 42 && Y == topY + 34) begin oled_data = 16'hffff; end
        else if (X == leftX + 43 && Y == topY + 34) begin oled_data = 16'h8f7d; end
        else if (X == leftX + 44 && Y == topY + 34) begin oled_data = 16'h2aca; end
        else if (X == leftX + 46 && Y == topY + 34) begin oled_data = 16'h2124; end
        else if (X == leftX + 48 && Y == topY + 34) begin oled_data = 16'h2945; end
        else if (X == leftX + 49 && Y == topY + 34) begin oled_data = 16'h31a6; end
        else if (X == leftX + 50 && Y == topY + 34) begin oled_data = 16'h39e7; end
        else if (X == leftX + 51 && Y == topY + 34) begin oled_data = 16'h29e7; end
        else if (X == leftX + 52 && Y == topY + 34) begin oled_data = 16'h21a5; end
        else if (X == leftX + 0 && Y == topY + 35) begin oled_data = 16'h2124; end
        else if (X == leftX + 8 && Y == topY + 35) begin oled_data = 16'h3166; end
        else if (X == leftX + 9 && Y == topY + 35) begin oled_data = 16'h72ac; end
        else if (X == leftX + 10 && Y == topY + 35) begin oled_data = 16'he6bb; end
        else if (X >= leftX + 11 && X <= leftX + 13 && Y == topY + 35) begin oled_data = 16'hffff; end
        else if (X == leftX + 14 && Y == topY + 35) begin oled_data = 16'heffd; end
        else if (X == leftX + 15 && Y == topY + 35) begin oled_data = 16'he7fc; end
        else if (X == leftX + 16 && Y == topY + 35) begin oled_data = 16'hf7fe; end
        else if (X == leftX + 17 && Y == topY + 35) begin oled_data = 16'hffff; end
        else if (X == leftX + 18 && Y == topY + 35) begin oled_data = 16'heffe; end
        else if (X == leftX + 19 && Y == topY + 35) begin oled_data = 16'h879b; end
        else if (X == leftX + 20 && Y == topY + 35) begin oled_data = 16'h2cd2; end
        else if (X == leftX + 21 && Y == topY + 35) begin oled_data = 16'h2185; end
        else if (X == leftX + 22 && Y == topY + 35) begin oled_data = 16'h29e5; end
        else if (X == leftX + 23 && Y == topY + 35) begin oled_data = 16'h33c6; end
        else if (X == leftX + 24 && Y == topY + 35) begin oled_data = 16'h33e5; end
        else if (X == leftX + 25 && Y == topY + 35) begin oled_data = 16'h33e5; end
        else if (X == leftX + 26 && Y == topY + 35) begin oled_data = 16'h4407; end
        else if (X == leftX + 27 && Y == topY + 35) begin oled_data = 16'hbb53; end
        else if (X == leftX + 28 && Y == topY + 35) begin oled_data = 16'hff7f; end
        else if (X == leftX + 29 && Y == topY + 35) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 35) begin oled_data = 16'hefff; end
        else if (X == leftX + 31 && Y == topY + 35) begin oled_data = 16'h3679; end
        else if (X == leftX + 32 && Y == topY + 35) begin oled_data = 16'h32c9; end
        else if (X == leftX + 33 && Y == topY + 35) begin oled_data = 16'hab53; end
        else if (X == leftX + 34 && Y == topY + 35) begin oled_data = 16'hff3f; end
        else if (X == leftX + 35 && Y == topY + 35) begin oled_data = 16'hffff; end
        else if (X == leftX + 36 && Y == topY + 35) begin oled_data = 16'hdfbe; end
        else if (X == leftX + 37 && Y == topY + 35) begin oled_data = 16'h3d95; end
        else if (X == leftX + 38 && Y == topY + 35) begin oled_data = 16'h2a08; end
        else if (X == leftX + 39 && Y == topY + 35) begin oled_data = 16'h59a9; end
        else if (X == leftX + 40 && Y == topY + 35) begin oled_data = 16'hdb18; end
        else if (X == leftX + 41 && Y == topY + 35) begin oled_data = 16'hffdf; end
        else if (X == leftX + 42 && Y == topY + 35) begin oled_data = 16'hffff; end
        else if (X == leftX + 43 && Y == topY + 35) begin oled_data = 16'hcfdf; end
        else if (X == leftX + 44 && Y == topY + 35) begin oled_data = 16'h3491; end
        else if (X == leftX + 45 && Y == topY + 35) begin oled_data = 16'h2965; end
        else if (X == leftX + 46 && Y == topY + 35) begin oled_data = 16'h5169; end
        else if (X == leftX + 47 && Y == topY + 35) begin oled_data = 16'ha353; end
        else if (X == leftX + 48 && Y == topY + 35) begin oled_data = 16'he65b; end
        else if (X == leftX + 49 && Y == topY + 35) begin oled_data = 16'hf7be; end
        else if (X == leftX + 50 && Y == topY + 35) begin oled_data = 16'hffff; end
        else if (X == leftX + 51 && Y == topY + 35) begin oled_data = 16'hf7df; end
        else if (X == leftX + 52 && Y == topY + 35) begin oled_data = 16'hc77d; end
        else if (X == leftX + 53 && Y == topY + 35) begin oled_data = 16'h5617; end
        else if (X == leftX + 54 && Y == topY + 35) begin oled_data = 16'h22cb; end
        else if (X == leftX + 0 && Y == topY + 36) begin oled_data = 16'h2124; end
        else if (X == leftX + 8 && Y == topY + 36) begin oled_data = 16'h3967; end
        else if (X == leftX + 9 && Y == topY + 36) begin oled_data = 16'h924f; end
        else if (X == leftX + 10 && Y == topY + 36) begin oled_data = 16'hfefe; end
        else if (X >= leftX + 11 && X <= leftX + 12 && Y == topY + 36) begin oled_data = 16'hffff; end
        else if (X == leftX + 13 && Y == topY + 36) begin oled_data = 16'h97f2; end
        else if (X == leftX + 14 && Y == topY + 36) begin oled_data = 16'h4648; end
        else if (X == leftX + 15 && Y == topY + 36) begin oled_data = 16'h5508; end
        else if (X == leftX + 16 && Y == topY + 36) begin oled_data = 16'hce37; end
        else if (X >= leftX + 17 && X <= leftX + 18 && Y == topY + 36) begin oled_data = 16'hffff; end
        else if (X == leftX + 19 && Y == topY + 36) begin oled_data = 16'h9ff7; end
        else if (X == leftX + 20 && Y == topY + 36) begin oled_data = 16'h2df5; end
        else if (X == leftX + 21 && Y == topY + 36) begin oled_data = 16'h2186; end
        else if (X == leftX + 26 && Y == topY + 36) begin oled_data = 16'h4167; end
        else if (X == leftX + 27 && Y == topY + 36) begin oled_data = 16'hc1f5; end
        else if (X == leftX + 28 && Y == topY + 36) begin oled_data = 16'hff7f; end
        else if (X == leftX + 29 && Y == topY + 36) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 36) begin oled_data = 16'hefff; end
        else if (X == leftX + 31 && Y == topY + 36) begin oled_data = 16'h3679; end
        else if (X == leftX + 32 && Y == topY + 36) begin oled_data = 16'h2a28; end
        else if (X == leftX + 33 && Y == topY + 36) begin oled_data = 16'h598a; end
        else if (X == leftX + 34 && Y == topY + 36) begin oled_data = 16'hed3b; end
        else if (X >= leftX + 35 && X <= leftX + 36 && Y == topY + 36) begin oled_data = 16'hffff; end
        else if (X == leftX + 37 && Y == topY + 36) begin oled_data = 16'h673c; end
        else if (X == leftX + 38 && Y == topY + 36) begin oled_data = 16'h3aec; end
        else if (X == leftX + 39 && Y == topY + 36) begin oled_data = 16'h79cd; end
        else if (X == leftX + 40 && Y == topY + 36) begin oled_data = 16'hf45c; end
        else if (X >= leftX + 41 && X <= leftX + 42 && Y == topY + 36) begin oled_data = 16'hffff; end
        else if (X == leftX + 43 && Y == topY + 36) begin oled_data = 16'h97be; end
        else if (X == leftX + 44 && Y == topY + 36) begin oled_data = 16'h2b0b; end
        else if (X == leftX + 45 && Y == topY + 36) begin oled_data = 16'h4187; end
        else if (X == leftX + 46 && Y == topY + 36) begin oled_data = 16'hb273; end
        else if (X == leftX + 47 && Y == topY + 36) begin oled_data = 16'hff5f; end
        else if (X >= leftX + 48 && X <= leftX + 52 && Y == topY + 36) begin oled_data = 16'hffff; end
        else if (X == leftX + 53 && Y == topY + 36) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 54 && Y == topY + 36) begin oled_data = 16'ha79e; end
        else if (X == leftX + 55 && Y == topY + 36) begin oled_data = 16'h4534; end
        else if (X == leftX + 56 && Y == topY + 36) begin oled_data = 16'h2289; end
        else if (X == leftX + 0 && Y == topY + 37) begin oled_data = 16'h2124; end
        else if (X == leftX + 8 && Y == topY + 37) begin oled_data = 16'h39a7; end
        else if (X == leftX + 9 && Y == topY + 37) begin oled_data = 16'h9ab0; end
        else if (X == leftX + 10 && Y == topY + 37) begin oled_data = 16'hff5f; end
        else if (X == leftX + 11 && Y == topY + 37) begin oled_data = 16'hffff; end
        else if (X == leftX + 12 && Y == topY + 37) begin oled_data = 16'hfffe; end
        else if (X == leftX + 13 && Y == topY + 37) begin oled_data = 16'h47d2; end
        else if (X == leftX + 14 && Y == topY + 37) begin oled_data = 16'h334c; end
        else if (X == leftX + 15 && Y == topY + 37) begin oled_data = 16'h5a6a; end
        else if (X == leftX + 16 && Y == topY + 37) begin oled_data = 16'hecbb; end
        else if (X >= leftX + 17 && X <= leftX + 18 && Y == topY + 37) begin oled_data = 16'hffff; end
        else if (X == leftX + 19 && Y == topY + 37) begin oled_data = 16'ha7f7; end
        else if (X == leftX + 20 && Y == topY + 37) begin oled_data = 16'h2e15; end
        else if (X == leftX + 21 && Y == topY + 37) begin oled_data = 16'h31a7; end
        else if (X == leftX + 22 && Y == topY + 37) begin oled_data = 16'h718c; end
        else if (X == leftX + 23 && Y == topY + 37) begin oled_data = 16'hb434; end
        else if (X == leftX + 24 && Y == topY + 37) begin oled_data = 16'hb5b6; end
        else if (X == leftX + 25 && Y == topY + 37) begin oled_data = 16'hb5b6; end
        else if (X == leftX + 26 && Y == topY + 37) begin oled_data = 16'hbdd7; end
        else if (X == leftX + 27 && Y == topY + 37) begin oled_data = 16'he61b; end
        else if (X == leftX + 28 && Y == topY + 37) begin oled_data = 16'hffdf; end
        else if (X == leftX + 29 && Y == topY + 37) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 37) begin oled_data = 16'he7ff; end
        else if (X == leftX + 31 && Y == topY + 37) begin oled_data = 16'h3e79; end
        else if (X == leftX + 32 && Y == topY + 37) begin oled_data = 16'h2a28; end
        else if (X == leftX + 33 && Y == topY + 37) begin oled_data = 16'h3967; end
        else if (X == leftX + 34 && Y == topY + 37) begin oled_data = 16'hc2f5; end
        else if (X >= leftX + 35 && X <= leftX + 36 && Y == topY + 37) begin oled_data = 16'hffff; end
        else if (X == leftX + 37 && Y == topY + 37) begin oled_data = 16'ha7df; end
        else if (X == leftX + 38 && Y == topY + 37) begin oled_data = 16'h4c52; end
        else if (X == leftX + 39 && Y == topY + 37) begin oled_data = 16'haa13; end
        else if (X == leftX + 40 && Y == topY + 37) begin oled_data = 16'hfe3e; end
        else if (X == leftX + 41 && Y == topY + 37) begin oled_data = 16'hffff; end
        else if (X == leftX + 42 && Y == topY + 37) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 43 && Y == topY + 37) begin oled_data = 16'h5679; end
        else if (X == leftX + 44 && Y == topY + 37) begin oled_data = 16'h2a07; end
        else if (X == leftX + 45 && Y == topY + 37) begin oled_data = 16'h59aa; end
        else if (X == leftX + 46 && Y == topY + 37) begin oled_data = 16'he3f9; end
        else if (X >= leftX + 47 && X <= leftX + 48 && Y == topY + 37) begin oled_data = 16'hffff; end
        else if (X == leftX + 49 && Y == topY + 37) begin oled_data = 16'hdfff; end
        else if (X == leftX + 50 && Y == topY + 37) begin oled_data = 16'h6fb9; end
        else if (X == leftX + 51 && Y == topY + 37) begin oled_data = 16'h8610; end
        else if (X == leftX + 52 && Y == topY + 37) begin oled_data = 16'hed7b; end
        else if (X >= leftX + 53 && X <= leftX + 54 && Y == topY + 37) begin oled_data = 16'hffff; end
        else if (X == leftX + 55 && Y == topY + 37) begin oled_data = 16'hcfff; end
        else if (X == leftX + 56 && Y == topY + 37) begin oled_data = 16'h2eba; end
        else if (X == leftX + 57 && Y == topY + 37) begin oled_data = 16'h21c6; end
        else if (X == leftX + 0 && Y == topY + 38) begin oled_data = 16'h2124; end
        else if (X == leftX + 8 && Y == topY + 38) begin oled_data = 16'h3186; end
        else if (X == leftX + 9 && Y == topY + 38) begin oled_data = 16'h6acb; end
        else if (X == leftX + 10 && Y == topY + 38) begin oled_data = 16'hee9c; end
        else if (X >= leftX + 11 && X <= leftX + 12 && Y == topY + 38) begin oled_data = 16'hffff; end
        else if (X == leftX + 13 && Y == topY + 38) begin oled_data = 16'h8fdc; end
        else if (X == leftX + 14 && Y == topY + 38) begin oled_data = 16'h3555; end
        else if (X == leftX + 15 && Y == topY + 38) begin oled_data = 16'h5aab; end
        else if (X == leftX + 16 && Y == topY + 38) begin oled_data = 16'hecdb; end
        else if (X >= leftX + 17 && X <= leftX + 18 && Y == topY + 38) begin oled_data = 16'hffff; end
        else if (X == leftX + 19 && Y == topY + 38) begin oled_data = 16'ha7f7; end
        else if (X == leftX + 20 && Y == topY + 38) begin oled_data = 16'h3616; end
        else if (X == leftX + 21 && Y == topY + 38) begin oled_data = 16'h6a0d; end
        else if (X == leftX + 22 && Y == topY + 38) begin oled_data = 16'hec3b; end
        else if (X == leftX + 23 && Y == topY + 38) begin oled_data = 16'hffbf; end
        else if (X >= leftX + 24 && X <= leftX + 29 && Y == topY + 38) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 38) begin oled_data = 16'h679d; end
        else if (X == leftX + 31 && Y == topY + 38) begin oled_data = 16'h336b; end
        else if (X == leftX + 32 && Y == topY + 38) begin oled_data = 16'h2165; end
        else if (X == leftX + 33 && Y == topY + 38) begin oled_data = 16'h4968; end
        else if (X == leftX + 34 && Y == topY + 38) begin oled_data = 16'hd2d7; end
        else if (X == leftX + 35 && Y == topY + 38) begin oled_data = 16'hff7f; end
        else if (X == leftX + 36 && Y == topY + 38) begin oled_data = 16'hffff; end
        else if (X == leftX + 37 && Y == topY + 38) begin oled_data = 16'hb7bf; end
        else if (X == leftX + 38 && Y == topY + 38) begin oled_data = 16'h94ba; end
        else if (X == leftX + 39 && Y == topY + 38) begin oled_data = 16'hec3b; end
        else if (X == leftX + 40 && Y == topY + 38) begin oled_data = 16'hffbf; end
        else if (X == leftX + 41 && Y == topY + 38) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 42 && Y == topY + 38) begin oled_data = 16'h9f9c; end
        else if (X == leftX + 43 && Y == topY + 38) begin oled_data = 16'h340e; end
        else if (X == leftX + 44 && Y == topY + 38) begin oled_data = 16'h3187; end
        else if (X == leftX + 45 && Y == topY + 38) begin oled_data = 16'h99f0; end
        else if (X == leftX + 46 && Y == topY + 38) begin oled_data = 16'hfebe; end
        else if (X == leftX + 47 && Y == topY + 38) begin oled_data = 16'hffff; end
        else if (X == leftX + 48 && Y == topY + 38) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 49 && Y == topY + 38) begin oled_data = 16'h57df; end
        else if (X == leftX + 50 && Y == topY + 38) begin oled_data = 16'h2b8d; end
        else if (X == leftX + 51 && Y == topY + 38) begin oled_data = 16'h3165; end
        else if (X == leftX + 52 && Y == topY + 38) begin oled_data = 16'h81ee; end
        else if (X == leftX + 53 && Y == topY + 38) begin oled_data = 16'hfdbd; end
        else if (X == leftX + 54 && Y == topY + 38) begin oled_data = 16'hefff; end
        else if (X == leftX + 55 && Y == topY + 38) begin oled_data = 16'hcfff; end
        else if (X == leftX + 56 && Y == topY + 38) begin oled_data = 16'h4fff; end
        else if (X == leftX + 57 && Y == topY + 38) begin oled_data = 16'h23ce; end
        else if (X == leftX + 59 && Y == topY + 38) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 39) begin oled_data = 16'h2124; end
        else if (X == leftX + 7 && Y == topY + 39) begin oled_data = 16'h2124; end
        else if (X == leftX + 8 && Y == topY + 39) begin oled_data = 16'h3166; end
        else if (X == leftX + 9 && Y == topY + 39) begin oled_data = 16'h6a8b; end
        else if (X == leftX + 10 && Y == topY + 39) begin oled_data = 16'hceb8; end
        else if (X >= leftX + 11 && X <= leftX + 13 && Y == topY + 39) begin oled_data = 16'hffff; end
        else if (X == leftX + 14 && Y == topY + 39) begin oled_data = 16'hdfdf; end
        else if (X == leftX + 15 && Y == topY + 39) begin oled_data = 16'hdf1c; end
        else if (X == leftX + 16 && Y == topY + 39) begin oled_data = 16'hf77e; end
        else if (X == leftX + 17 && Y == topY + 39) begin oled_data = 16'hffff; end
        else if (X == leftX + 18 && Y == topY + 39) begin oled_data = 16'hcff9; end
        else if (X == leftX + 19 && Y == topY + 39) begin oled_data = 16'h4f6d; end
        else if (X == leftX + 20 && Y == topY + 39) begin oled_data = 16'h3329; end
        else if (X == leftX + 21 && Y == topY + 39) begin oled_data = 16'h51e9; end
        else if (X == leftX + 22 && Y == topY + 39) begin oled_data = 16'had13; end
        else if (X == leftX + 23 && Y == topY + 39) begin oled_data = 16'haff5; end
        else if (X == leftX + 24 && Y == topY + 39) begin oled_data = 16'haff5; end
        else if (X == leftX + 25 && Y == topY + 39) begin oled_data = 16'haff5; end
        else if (X == leftX + 26 && Y == topY + 39) begin oled_data = 16'hcf58; end
        else if (X == leftX + 27 && Y == topY + 39) begin oled_data = 16'hff7f; end
        else if (X >= leftX + 28 && X <= leftX + 29 && Y == topY + 39) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 39) begin oled_data = 16'h4f3c; end
        else if (X == leftX + 31 && Y == topY + 39) begin oled_data = 16'h2a89; end
        else if (X == leftX + 33 && Y == topY + 39) begin oled_data = 16'h3967; end
        else if (X == leftX + 34 && Y == topY + 39) begin oled_data = 16'hcb35; end
        else if (X >= leftX + 35 && X <= leftX + 36 && Y == topY + 39) begin oled_data = 16'hffff; end
        else if (X == leftX + 37 && Y == topY + 39) begin oled_data = 16'h97bf; end
        else if (X == leftX + 38 && Y == topY + 39) begin oled_data = 16'hcc1c; end
        else if (X == leftX + 39 && Y == topY + 39) begin oled_data = 16'hffdf; end
        else if (X == leftX + 40 && Y == topY + 39) begin oled_data = 16'hffff; end
        else if (X == leftX + 41 && Y == topY + 39) begin oled_data = 16'hb7ff; end
        else if (X == leftX + 42 && Y == topY + 39) begin oled_data = 16'h3490; end
        else if (X == leftX + 43 && Y == topY + 39) begin oled_data = 16'h2185; end
        else if (X == leftX + 44 && Y == topY + 39) begin oled_data = 16'h4188; end
        else if (X == leftX + 45 && Y == topY + 39) begin oled_data = 16'hc235; end
        else if (X == leftX + 46 && Y == topY + 39) begin oled_data = 16'he75f; end
        else if (X == leftX + 47 && Y == topY + 39) begin oled_data = 16'hd7ff; end
        else if (X == leftX + 48 && Y == topY + 39) begin oled_data = 16'hafff; end
        else if (X == leftX + 49 && Y == topY + 39) begin oled_data = 16'h2eba; end
        else if (X == leftX + 50 && Y == topY + 39) begin oled_data = 16'h21a6; end
        else if (X == leftX + 52 && Y == topY + 39) begin oled_data = 16'h51a9; end
        else if (X == leftX + 53 && Y == topY + 39) begin oled_data = 16'hdb18; end
        else if (X == leftX + 54 && Y == topY + 39) begin oled_data = 16'hcf7f; end
        else if (X == leftX + 55 && Y == topY + 39) begin oled_data = 16'h97df; end
        else if (X == leftX + 56 && Y == topY + 39) begin oled_data = 16'h7fff; end
        else if (X == leftX + 57 && Y == topY + 39) begin oled_data = 16'h2db6; end
        else if (X == leftX + 58 && Y == topY + 39) begin oled_data = 16'h2165; end
        else if (X == leftX + 0 && Y == topY + 40) begin oled_data = 16'h2124; end
        else if (X == leftX + 7 && Y == topY + 40) begin oled_data = 16'h2124; end
        else if (X == leftX + 9 && Y == topY + 40) begin oled_data = 16'h41e7; end
        else if (X == leftX + 10 && Y == topY + 40) begin oled_data = 16'h8c8f; end
        else if (X == leftX + 11 && Y == topY + 40) begin oled_data = 16'hefdc; end
        else if (X >= leftX + 12 && X <= leftX + 17 && Y == topY + 40) begin oled_data = 16'hffff; end
        else if (X == leftX + 18 && Y == topY + 40) begin oled_data = 16'hbff8; end
        else if (X == leftX + 19 && Y == topY + 40) begin oled_data = 16'h2ed6; end
        else if (X == leftX + 20 && Y == topY + 40) begin oled_data = 16'h21c6; end
        else if (X == leftX + 21 && Y == topY + 40) begin oled_data = 16'h2164; end
        else if (X == leftX + 22 && Y == topY + 40) begin oled_data = 16'h2a05; end
        else if (X == leftX + 23 && Y == topY + 40) begin oled_data = 16'h2a65; end
        else if (X == leftX + 24 && Y == topY + 40) begin oled_data = 16'h2a65; end
        else if (X == leftX + 25 && Y == topY + 40) begin oled_data = 16'h3265; end
        else if (X == leftX + 26 && Y == topY + 40) begin oled_data = 16'h7aad; end
        else if (X == leftX + 27 && Y == topY + 40) begin oled_data = 16'he55a; end
        else if (X == leftX + 28 && Y == topY + 40) begin oled_data = 16'hffbf; end
        else if (X == leftX + 29 && Y == topY + 40) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 40) begin oled_data = 16'h9f7d; end
        else if (X == leftX + 31 && Y == topY + 40) begin oled_data = 16'h2c50; end
        else if (X == leftX + 32 && Y == topY + 40) begin oled_data = 16'h21a6; end
        else if (X == leftX + 33 && Y == topY + 40) begin oled_data = 16'h2945; end
        else if (X == leftX + 34 && Y == topY + 40) begin oled_data = 16'h720c; end
        else if (X == leftX + 35 && Y == topY + 40) begin oled_data = 16'heedc; end
        else if (X == leftX + 36 && Y == topY + 40) begin oled_data = 16'hffdf; end
        else if (X == leftX + 37 && Y == topY + 40) begin oled_data = 16'hcfff; end
        else if (X == leftX + 38 && Y == topY + 40) begin oled_data = 16'haf3e; end
        else if (X == leftX + 39 && Y == topY + 40) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 40 && Y == topY + 40) begin oled_data = 16'hffff; end
        else if (X == leftX + 41 && Y == topY + 40) begin oled_data = 16'h8f7d; end
        else if (X == leftX + 42 && Y == topY + 40) begin oled_data = 16'h2b0b; end
        else if (X == leftX + 43 && Y == topY + 40) begin oled_data = 16'h3166; end
        else if (X == leftX + 44 && Y == topY + 40) begin oled_data = 16'h81ce; end
        else if (X == leftX + 45 && Y == topY + 40) begin oled_data = 16'he4ba; end
        else if (X == leftX + 46 && Y == topY + 40) begin oled_data = 16'hbf1e; end
        else if (X == leftX + 47 && Y == topY + 40) begin oled_data = 16'h87df; end
        else if (X == leftX + 48 && Y == topY + 40) begin oled_data = 16'h37dd; end
        else if (X == leftX + 49 && Y == topY + 40) begin oled_data = 16'h2c6f; end
        else if (X == leftX + 51 && Y == topY + 40) begin oled_data = 16'h2945; end
        else if (X == leftX + 52 && Y == topY + 40) begin oled_data = 16'h69ac; end
        else if (X == leftX + 53 && Y == topY + 40) begin oled_data = 16'hdc19; end
        else if (X == leftX + 54 && Y == topY + 40) begin oled_data = 16'hcebe; end
        else if (X == leftX + 55 && Y == topY + 40) begin oled_data = 16'hb7df; end
        else if (X == leftX + 56 && Y == topY + 40) begin oled_data = 16'h7fff; end
        else if (X == leftX + 57 && Y == topY + 40) begin oled_data = 16'h34f2; end
        else if (X == leftX + 58 && Y == topY + 40) begin oled_data = 16'h2164; end
        else if (X == leftX + 0 && Y == topY + 41) begin oled_data = 16'h2124; end
        else if (X == leftX + 8 && Y == topY + 41) begin oled_data = 16'h2945; end
        else if (X == leftX + 9 && Y == topY + 41) begin oled_data = 16'h6a2b; end
        else if (X == leftX + 10 && Y == topY + 41) begin oled_data = 16'hcdf8; end
        else if (X >= leftX + 11 && X <= leftX + 12 && Y == topY + 41) begin oled_data = 16'hffff; end
        else if (X == leftX + 13 && Y == topY + 41) begin oled_data = 16'heffd; end
        else if (X == leftX + 14 && Y == topY + 41) begin oled_data = 16'h77f2; end
        else if (X == leftX + 15 && Y == topY + 41) begin oled_data = 16'h8fb1; end
        else if (X == leftX + 16 && Y == topY + 41) begin oled_data = 16'he7fb; end
        else if (X == leftX + 17 && Y == topY + 41) begin oled_data = 16'hffff; end
        else if (X == leftX + 18 && Y == topY + 41) begin oled_data = 16'hd7fb; end
        else if (X == leftX + 19 && Y == topY + 41) begin oled_data = 16'h5719; end
        else if (X == leftX + 20 && Y == topY + 41) begin oled_data = 16'h232c; end
        else if (X == leftX + 21 && Y == topY + 41) begin oled_data = 16'h2145; end
        else if (X == leftX + 25 && Y == topY + 41) begin oled_data = 16'h2944; end
        else if (X == leftX + 26 && Y == topY + 41) begin oled_data = 16'h598a; end
        else if (X == leftX + 27 && Y == topY + 41) begin oled_data = 16'hd337; end
        else if (X == leftX + 28 && Y == topY + 41) begin oled_data = 16'hff9f; end
        else if (X == leftX + 29 && Y == topY + 41) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 41) begin oled_data = 16'hcfff; end
        else if (X == leftX + 31 && Y == topY + 41) begin oled_data = 16'h3dd6; end
        else if (X == leftX + 32 && Y == topY + 41) begin oled_data = 16'h29e7; end
        else if (X == leftX + 34 && Y == topY + 41) begin oled_data = 16'h39a6; end
        else if (X == leftX + 35 && Y == topY + 41) begin oled_data = 16'hb293; end
        else if (X == leftX + 36 && Y == topY + 41) begin oled_data = 16'hfe5e; end
        else if (X == leftX + 37 && Y == topY + 41) begin oled_data = 16'hffff; end
        else if (X == leftX + 38 && Y == topY + 41) begin oled_data = 16'hd7ff; end
        else if (X == leftX + 39 && Y == topY + 41) begin oled_data = 16'he7ff; end
        else if (X == leftX + 40 && Y == topY + 41) begin oled_data = 16'hffff; end
        else if (X == leftX + 41 && Y == topY + 41) begin oled_data = 16'hbfde; end
        else if (X == leftX + 42 && Y == topY + 41) begin oled_data = 16'h3450; end
        else if (X == leftX + 43 && Y == topY + 41) begin oled_data = 16'h41a7; end
        else if (X == leftX + 44 && Y == topY + 41) begin oled_data = 16'hb9f4; end
        else if (X == leftX + 45 && Y == topY + 41) begin oled_data = 16'hd63e; end
        else if (X == leftX + 46 && Y == topY + 41) begin oled_data = 16'h8fdf; end
        else if (X == leftX + 47 && Y == topY + 41) begin oled_data = 16'h6fff; end
        else if (X == leftX + 48 && Y == topY + 41) begin oled_data = 16'h2f1b; end
        else if (X == leftX + 49 && Y == topY + 41) begin oled_data = 16'h21c6; end
        else if (X == leftX + 50 && Y == topY + 41) begin oled_data = 16'h2124; end
        else if (X == leftX + 51 && Y == topY + 41) begin oled_data = 16'h3165; end
        else if (X == leftX + 52 && Y == topY + 41) begin oled_data = 16'h91d0; end
        else if (X == leftX + 53 && Y == topY + 41) begin oled_data = 16'hf57d; end
        else if (X == leftX + 54 && Y == topY + 41) begin oled_data = 16'hdfdf; end
        else if (X == leftX + 55 && Y == topY + 41) begin oled_data = 16'hf7ff; end
        else if (X == leftX + 56 && Y == topY + 41) begin oled_data = 16'h3fbe; end
        else if (X == leftX + 57 && Y == topY + 41) begin oled_data = 16'h2289; end
        else if (X == leftX + 0 && Y == topY + 42) begin oled_data = 16'h2124; end
        else if (X == leftX + 8 && Y == topY + 42) begin oled_data = 16'h3145; end
        else if (X == leftX + 9 && Y == topY + 42) begin oled_data = 16'h6a4b; end
        else if (X == leftX + 10 && Y == topY + 42) begin oled_data = 16'hcd57; end
        else if (X == leftX + 11 && Y == topY + 42) begin oled_data = 16'hffff; end
        else if (X == leftX + 12 && Y == topY + 42) begin oled_data = 16'hf7fe; end
        else if (X == leftX + 13 && Y == topY + 42) begin oled_data = 16'hbff7; end
        else if (X == leftX + 14 && Y == topY + 42) begin oled_data = 16'h46d1; end
        else if (X == leftX + 15 && Y == topY + 42) begin oled_data = 16'h6bce; end
        else if (X == leftX + 16 && Y == topY + 42) begin oled_data = 16'hde19; end
        else if (X == leftX + 17 && Y == topY + 42) begin oled_data = 16'hffff; end
        else if (X == leftX + 18 && Y == topY + 42) begin oled_data = 16'hf7fe; end
        else if (X == leftX + 19 && Y == topY + 42) begin oled_data = 16'h97f6; end
        else if (X == leftX + 20 && Y == topY + 42) begin oled_data = 16'h3594; end
        else if (X == leftX + 21 && Y == topY + 42) begin oled_data = 16'h59cb; end
        else if (X == leftX + 22 && Y == topY + 42) begin oled_data = 16'h9351; end
        else if (X == leftX + 23 && Y == topY + 42) begin oled_data = 16'h9cd2; end
        else if (X == leftX + 24 && Y == topY + 42) begin oled_data = 16'h94d2; end
        else if (X == leftX + 25 && Y == topY + 42) begin oled_data = 16'h9cf3; end
        else if (X == leftX + 26 && Y == topY + 42) begin oled_data = 16'hd539; end
        else if (X == leftX + 27 && Y == topY + 42) begin oled_data = 16'hff5f; end
        else if (X >= leftX + 28 && X <= leftX + 29 && Y == topY + 42) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 42) begin oled_data = 16'h879d; end
        else if (X == leftX + 31 && Y == topY + 42) begin oled_data = 16'h3490; end
        else if (X == leftX + 32 && Y == topY + 42) begin oled_data = 16'h21a5; end
        else if (X == leftX + 34 && Y == topY + 42) begin oled_data = 16'h3165; end
        else if (X == leftX + 35 && Y == topY + 42) begin oled_data = 16'h8b0f; end
        else if (X == leftX + 36 && Y == topY + 42) begin oled_data = 16'hf71e; end
        else if (X >= leftX + 37 && X <= leftX + 39 && Y == topY + 42) begin oled_data = 16'hffff; end
        else if (X == leftX + 40 && Y == topY + 42) begin oled_data = 16'hcfff; end
        else if (X == leftX + 41 && Y == topY + 42) begin oled_data = 16'h45d4; end
        else if (X == leftX + 42 && Y == topY + 42) begin oled_data = 16'h29e6; end
        else if (X == leftX + 43 && Y == topY + 42) begin oled_data = 16'h3166; end
        else if (X == leftX + 44 && Y == topY + 42) begin oled_data = 16'ha1f1; end
        else if (X == leftX + 45 && Y == topY + 42) begin oled_data = 16'hfefe; end
        else if (X == leftX + 46 && Y == topY + 42) begin oled_data = 16'hffff; end
        else if (X == leftX + 47 && Y == topY + 42) begin oled_data = 16'hdfff; end
        else if (X == leftX + 48 && Y == topY + 42) begin oled_data = 16'h3f5c; end
        else if (X == leftX + 49 && Y == topY + 42) begin oled_data = 16'h2228; end
        else if (X == leftX + 51 && Y == topY + 42) begin oled_data = 16'h3166; end
        else if (X == leftX + 52 && Y == topY + 42) begin oled_data = 16'h99f1; end
        else if (X == leftX + 53 && Y == topY + 42) begin oled_data = 16'hf69e; end
        else if (X == leftX + 54 && Y == topY + 42) begin oled_data = 16'hefff; end
        else if (X == leftX + 55 && Y == topY + 42) begin oled_data = 16'hdfff; end
        else if (X == leftX + 56 && Y == topY + 42) begin oled_data = 16'h3f9d; end
        else if (X == leftX + 57 && Y == topY + 42) begin oled_data = 16'h2268; end
        else if (X == leftX + 0 && Y == topY + 43) begin oled_data = 16'h2124; end
        else if (X == leftX + 6 && Y == topY + 43) begin oled_data = 16'h2124; end
        else if (X == leftX + 7 && Y == topY + 43) begin oled_data = 16'h2945; end
        else if (X == leftX + 8 && Y == topY + 43) begin oled_data = 16'h5a09; end
        else if (X == leftX + 9 && Y == topY + 43) begin oled_data = 16'hc516; end
        else if (X == leftX + 10 && Y == topY + 43) begin oled_data = 16'hf7fe; end
        else if (X == leftX + 11 && Y == topY + 43) begin oled_data = 16'hffff; end
        else if (X == leftX + 12 && Y == topY + 43) begin oled_data = 16'hc7d9; end
        else if (X == leftX + 13 && Y == topY + 43) begin oled_data = 16'h4771; end
        else if (X == leftX + 14 && Y == topY + 43) begin oled_data = 16'h4bed; end
        else if (X == leftX + 15 && Y == topY + 43) begin oled_data = 16'hbc34; end
        else if (X == leftX + 16 && Y == topY + 43) begin oled_data = 16'he7fc; end
        else if (X == leftX + 17 && Y == topY + 43) begin oled_data = 16'hffff; end
        else if (X == leftX + 18 && Y == topY + 43) begin oled_data = 16'hd7fa; end
        else if (X == leftX + 19 && Y == topY + 43) begin oled_data = 16'h4f52; end
        else if (X == leftX + 20 && Y == topY + 43) begin oled_data = 16'h2b2a; end
        else if (X == leftX + 21 && Y == topY + 43) begin oled_data = 16'h61ab; end
        else if (X == leftX + 22 && Y == topY + 43) begin oled_data = 16'he399; end
        else if (X >= leftX + 23 && X <= leftX + 29 && Y == topY + 43) begin oled_data = 16'hffff; end
        else if (X == leftX + 30 && Y == topY + 43) begin oled_data = 16'hd7ff; end
        else if (X == leftX + 31 && Y == topY + 43) begin oled_data = 16'h3e37; end
        else if (X == leftX + 32 && Y == topY + 43) begin oled_data = 16'h2a07; end
        else if (X == leftX + 33 && Y == topY + 43) begin oled_data = 16'h2124; end
        else if (X == leftX + 35 && Y == topY + 43) begin oled_data = 16'h51e9; end
        else if (X == leftX + 36 && Y == topY + 43) begin oled_data = 16'hdaf7; end
        else if (X == leftX + 37 && Y == topY + 43) begin oled_data = 16'hff9f; end
        else if (X >= leftX + 38 && X <= leftX + 39 && Y == topY + 43) begin oled_data = 16'hffff; end
        else if (X == leftX + 40 && Y == topY + 43) begin oled_data = 16'hdfff; end
        else if (X == leftX + 41 && Y == topY + 43) begin oled_data = 16'h45d6; end
        else if (X == leftX + 42 && Y == topY + 43) begin oled_data = 16'h29e7; end
        else if (X == leftX + 44 && Y == topY + 43) begin oled_data = 16'h49a8; end
        else if (X == leftX + 45 && Y == topY + 43) begin oled_data = 16'hbad4; end
        else if (X == leftX + 46 && Y == topY + 43) begin oled_data = 16'hff5f; end
        else if (X == leftX + 47 && Y == topY + 43) begin oled_data = 16'hffff; end
        else if (X == leftX + 48 && Y == topY + 43) begin oled_data = 16'hdfdf; end
        else if (X == leftX + 49 && Y == topY + 43) begin oled_data = 16'h36fb; end
        else if (X == leftX + 50 && Y == topY + 43) begin oled_data = 16'h2207; end
        else if (X == leftX + 51 && Y == topY + 43) begin oled_data = 16'h2944; end
        else if (X == leftX + 52 && Y == topY + 43) begin oled_data = 16'h69ab; end
        else if (X == leftX + 53 && Y == topY + 43) begin oled_data = 16'hec5b; end
        else if (X >= leftX + 54 && X <= leftX + 55 && Y == topY + 43) begin oled_data = 16'hffff; end
        else if (X == leftX + 56 && Y == topY + 43) begin oled_data = 16'h8fff; end
        else if (X == leftX + 57 && Y == topY + 43) begin oled_data = 16'h2d13; end
        else if (X == leftX + 0 && Y == topY + 44) begin oled_data = 16'h2124; end
        else if (X == leftX + 8 && Y == topY + 44) begin oled_data = 16'h41a7; end
        else if (X == leftX + 9 && Y == topY + 44) begin oled_data = 16'h8bef; end
        else if (X == leftX + 10 && Y == topY + 44) begin oled_data = 16'hf7be; end
        else if (X == leftX + 11 && Y == topY + 44) begin oled_data = 16'hffff; end
        else if (X == leftX + 12 && Y == topY + 44) begin oled_data = 16'hf7fe; end
        else if (X == leftX + 13 && Y == topY + 44) begin oled_data = 16'h5fd5; end
        else if (X == leftX + 14 && Y == topY + 44) begin oled_data = 16'h3c2f; end
        else if (X == leftX + 15 && Y == topY + 44) begin oled_data = 16'h5b2a; end
        else if (X == leftX + 16 && Y == topY + 44) begin oled_data = 16'hce18; end
        else if (X >= leftX + 17 && X <= leftX + 18 && Y == topY + 44) begin oled_data = 16'hffff; end
        else if (X == leftX + 19 && Y == topY + 44) begin oled_data = 16'h9ff9; end
        else if (X == leftX + 20 && Y == topY + 44) begin oled_data = 16'h3df6; end
        else if (X == leftX + 21 && Y == topY + 44) begin oled_data = 16'h9af1; end
        else if (X == leftX + 22 && Y == topY + 44) begin oled_data = 16'hc798; end
        else if (X == leftX + 23 && Y == topY + 44) begin oled_data = 16'hc7f8; end
        else if (X == leftX + 24 && Y == topY + 44) begin oled_data = 16'hc7f8; end
        else if (X == leftX + 25 && Y == topY + 44) begin oled_data = 16'hc7f8; end
        else if (X == leftX + 26 && Y == topY + 44) begin oled_data = 16'hc7f8; end
        else if (X == leftX + 27 && Y == topY + 44) begin oled_data = 16'hc7f8; end
        else if (X == leftX + 28 && Y == topY + 44) begin oled_data = 16'hc7f8; end
        else if (X == leftX + 29 && Y == topY + 44) begin oled_data = 16'hc7f8; end
        else if (X == leftX + 30 && Y == topY + 44) begin oled_data = 16'h56b6; end
        else if (X == leftX + 31 && Y == topY + 44) begin oled_data = 16'h2ac9; end
        else if (X == leftX + 34 && Y == topY + 44) begin oled_data = 16'h2124; end
        else if (X == leftX + 35 && Y == topY + 44) begin oled_data = 16'h39a6; end
        else if (X == leftX + 36 && Y == topY + 44) begin oled_data = 16'h8510; end
        else if (X == leftX + 37 && Y == topY + 44) begin oled_data = 16'haff5; end
        else if (X == leftX + 38 && Y == topY + 44) begin oled_data = 16'hb7f5; end
        else if (X == leftX + 39 && Y == topY + 44) begin oled_data = 16'ha7b5; end
        else if (X == leftX + 40 && Y == topY + 44) begin oled_data = 16'h4572; end
        else if (X == leftX + 41 && Y == topY + 44) begin oled_data = 16'h2a26; end
        else if (X == leftX + 44 && Y == topY + 44) begin oled_data = 16'h4988; end
        else if (X == leftX + 45 && Y == topY + 44) begin oled_data = 16'hcb16; end
        else if (X == leftX + 46 && Y == topY + 44) begin oled_data = 16'hff9f; end
        else if (X == leftX + 47 && Y == topY + 44) begin oled_data = 16'hffff; end
        else if (X == leftX + 48 && Y == topY + 44) begin oled_data = 16'hdfff; end
        else if (X == leftX + 49 && Y == topY + 44) begin oled_data = 16'h473c; end
        else if (X == leftX + 50 && Y == topY + 44) begin oled_data = 16'h326a; end
        else if (X == leftX + 51 && Y == topY + 44) begin oled_data = 16'h79cd; end
        else if (X == leftX + 52 && Y == topY + 44) begin oled_data = 16'hd559; end
        else if (X == leftX + 53 && Y == topY + 44) begin oled_data = 16'hff7f; end
        else if (X == leftX + 54 && Y == topY + 44) begin oled_data = 16'hffff; end
        else if (X == leftX + 55 && Y == topY + 44) begin oled_data = 16'h9ffe; end
        else if (X == leftX + 56 && Y == topY + 44) begin oled_data = 16'h46b3; end
        else if (X == leftX + 57 && Y == topY + 44) begin oled_data = 16'h2a67; end
        else if (X == leftX + 58 && Y == topY + 44) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 45) begin oled_data = 16'h2124; end
        else if (X == leftX + 7 && Y == topY + 45) begin oled_data = 16'h41a7; end
        else if (X == leftX + 8 && Y == topY + 45) begin oled_data = 16'hb2f3; end
        else if (X == leftX + 9 && Y == topY + 45) begin oled_data = 16'hef9d; end
        else if (X == leftX + 10 && Y == topY + 45) begin oled_data = 16'hf7fe; end
        else if (X == leftX + 11 && Y == topY + 45) begin oled_data = 16'he7fc; end
        else if (X == leftX + 12 && Y == topY + 45) begin oled_data = 16'h4f8c; end
        else if (X == leftX + 13 && Y == topY + 45) begin oled_data = 16'h3467; end
        else if (X == leftX + 14 && Y == topY + 45) begin oled_data = 16'h5229; end
        else if (X == leftX + 15 && Y == topY + 45) begin oled_data = 16'hcbf6; end
        else if (X == leftX + 16 && Y == topY + 45) begin oled_data = 16'hefde; end
        else if (X == leftX + 17 && Y == topY + 45) begin oled_data = 16'hf7fe; end
        else if (X == leftX + 18 && Y == topY + 45) begin oled_data = 16'hbff7; end
        else if (X == leftX + 19 && Y == topY + 45) begin oled_data = 16'h3f0d; end
        else if (X == leftX + 20 && Y == topY + 45) begin oled_data = 16'h2a67; end
        else if (X == leftX + 21 && Y == topY + 45) begin oled_data = 16'h29e5; end
        else if (X == leftX + 22 && Y == topY + 45) begin oled_data = 16'h3325; end
        else if (X == leftX + 23 && Y == topY + 45) begin oled_data = 16'h2b45; end
        else if (X == leftX + 24 && Y == topY + 45) begin oled_data = 16'h2b25; end
        else if (X == leftX + 25 && Y == topY + 45) begin oled_data = 16'h2b25; end
        else if (X == leftX + 26 && Y == topY + 45) begin oled_data = 16'h2b45; end
        else if (X == leftX + 27 && Y == topY + 45) begin oled_data = 16'h2b45; end
        else if (X == leftX + 28 && Y == topY + 45) begin oled_data = 16'h2b45; end
        else if (X == leftX + 29 && Y == topY + 45) begin oled_data = 16'h3325; end
        else if (X == leftX + 30 && Y == topY + 45) begin oled_data = 16'h2a25; end
        else if (X == leftX + 34 && Y == topY + 45) begin oled_data = 16'h2124; end
        else if (X == leftX + 36 && Y == topY + 45) begin oled_data = 16'h29e5; end
        else if (X == leftX + 37 && Y == topY + 45) begin oled_data = 16'h2aa5; end
        else if (X == leftX + 38 && Y == topY + 45) begin oled_data = 16'h32a5; end
        else if (X == leftX + 39 && Y == topY + 45) begin oled_data = 16'h2a65; end
        else if (X == leftX + 40 && Y == topY + 45) begin oled_data = 16'h2184; end
        else if (X == leftX + 44 && Y == topY + 45) begin oled_data = 16'h2965; end
        else if (X == leftX + 45 && Y == topY + 45) begin oled_data = 16'h5a8a; end
        else if (X == leftX + 46 && Y == topY + 45) begin oled_data = 16'hc475; end
        else if (X == leftX + 47 && Y == topY + 45) begin oled_data = 16'hff3f; end
        else if (X == leftX + 48 && Y == topY + 45) begin oled_data = 16'hffff; end
        else if (X == leftX + 49 && Y == topY + 45) begin oled_data = 16'hefff; end
        else if (X == leftX + 50 && Y == topY + 45) begin oled_data = 16'hcf5d; end
        else if (X == leftX + 51 && Y == topY + 45) begin oled_data = 16'hdebd; end
        else if (X >= leftX + 52 && X <= leftX + 54 && Y == topY + 45) begin oled_data = 16'hffff; end
        else if (X == leftX + 55 && Y == topY + 45) begin oled_data = 16'h87ff; end
        else if (X == leftX + 56 && Y == topY + 45) begin oled_data = 16'h2cf3; end
        else if (X == leftX + 57 && Y == topY + 45) begin oled_data = 16'h2165; end
        else if (X == leftX + 0 && Y == topY + 46) begin oled_data = 16'h2124; end
        else if (X == leftX + 5 && Y == topY + 46) begin oled_data = 16'h2124; end
        else if (X == leftX + 7 && Y == topY + 46) begin oled_data = 16'h2184; end
        else if (X == leftX + 8 && Y == topY + 46) begin oled_data = 16'h3ac6; end
        else if (X == leftX + 9 && Y == topY + 46) begin oled_data = 16'h44e7; end
        else if (X == leftX + 10 && Y == topY + 46) begin oled_data = 16'h4507; end
        else if (X == leftX + 11 && Y == topY + 46) begin oled_data = 16'h3d07; end
        else if (X == leftX + 12 && Y == topY + 46) begin oled_data = 16'h2b26; end
        else if (X == leftX + 13 && Y == topY + 46) begin oled_data = 16'h2164; end
        else if (X == leftX + 14 && Y == topY + 46) begin oled_data = 16'h2985; end
        else if (X == leftX + 15 && Y == topY + 46) begin oled_data = 16'h3ae7; end
        else if (X == leftX + 16 && Y == topY + 46) begin oled_data = 16'h44e7; end
        else if (X == leftX + 17 && Y == topY + 46) begin oled_data = 16'h4507; end
        else if (X == leftX + 18 && Y == topY + 46) begin oled_data = 16'h3ce7; end
        else if (X == leftX + 19 && Y == topY + 46) begin oled_data = 16'h2aa6; end
        else if (X >= leftX + 43 && X <= leftX + 44 && Y == topY + 46) begin oled_data = 16'h2124; end
        else if (X == leftX + 45 && Y == topY + 46) begin oled_data = 16'h2945; end
        else if (X == leftX + 46 && Y == topY + 46) begin oled_data = 16'h69cb; end
        else if (X == leftX + 47 && Y == topY + 46) begin oled_data = 16'hecdb; end
        else if (X >= leftX + 48 && X <= leftX + 52 && Y == topY + 46) begin oled_data = 16'hffff; end
        else if (X == leftX + 53 && Y == topY + 46) begin oled_data = 16'hcfff; end
        else if (X == leftX + 54 && Y == topY + 46) begin oled_data = 16'h87d6; end
        else if (X == leftX + 55 && Y == topY + 46) begin oled_data = 16'h3e30; end
        else if (X == leftX + 56 && Y == topY + 46) begin oled_data = 16'h21c6; end
        else if (X == leftX + 0 && Y == topY + 47) begin oled_data = 16'h2124; end
        else if (X == leftX + 46 && Y == topY + 47) begin oled_data = 16'h2985; end
        else if (X == leftX + 47 && Y == topY + 47) begin oled_data = 16'h52e9; end
        else if (X == leftX + 48 && Y == topY + 47) begin oled_data = 16'h8dd0; end
        else if (X == leftX + 49 && Y == topY + 47) begin oled_data = 16'hb7b5; end
        else if (X == leftX + 50 && Y == topY + 47) begin oled_data = 16'hb7f6; end
        else if (X == leftX + 51 && Y == topY + 47) begin oled_data = 16'ha7f5; end
        else if (X == leftX + 52 && Y == topY + 47) begin oled_data = 16'h77b2; end
        else if (X == leftX + 53 && Y == topY + 47) begin oled_data = 16'h3dcc; end
        else if (X == leftX + 54 && Y == topY + 47) begin oled_data = 16'h2a66; end
        else if (X == leftX + 55 && Y == topY + 47) begin oled_data = 16'h2164; end
        else if (X == leftX + 57 && Y == topY + 47) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 48) begin oled_data = 16'h2124; end
        else if (X == leftX + 48 && Y == topY + 48) begin oled_data = 16'h2184; end
        else if (X == leftX + 49 && Y == topY + 48) begin oled_data = 16'h2a05; end
        else if (X == leftX + 50 && Y == topY + 48) begin oled_data = 16'h2a45; end
        else if (X == leftX + 51 && Y == topY + 48) begin oled_data = 16'h2a25; end
        else if (X == leftX + 52 && Y == topY + 48) begin oled_data = 16'h29c5; end
        else if (X == leftX + 54 && Y == topY + 48) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 49) begin oled_data = 16'h2124; end
        else if (X == leftX + 47 && Y == topY + 49) begin oled_data = 16'h2124; end
        else if (X == leftX + 54 && Y == topY + 49) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 50) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 51) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 52) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 53) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 54) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 55) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 56) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 57) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 58) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 59) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 60) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 61) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 62) begin oled_data = 16'h2124; end
        else if (X == leftX + 0 && Y == topY + 63) begin oled_data = 16'h2124; end
        else begin oled_data = 16'h2144; end
    end
endmodule
