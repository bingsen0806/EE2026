`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 24.03.2021 20:17:21
// Design Name: 
// Module Name: Stadium
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Stadium(
    input[6:0] X, 
    input [5:0] Y, 
    output reg [15:0] oled_data = 16'b0
    );
    always @ (X or Y) begin
    if (X == 0 && Y == 0) begin oled_data = 16'hce57; end
    else if (X == 1 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 2 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 3 && Y == 0) begin oled_data = 16'ha593; end
    else if (X == 4 && Y == 0) begin oled_data = 16'ha593; end
    else if (X == 5 && Y == 0) begin oled_data = 16'ha593; end
    else if (X == 6 && Y == 0) begin oled_data = 16'ha593; end
    else if (X == 7 && Y == 0) begin oled_data = 16'ha593; end
    else if (X == 8 && Y == 0) begin oled_data = 16'ha593; end
    else if (X == 9 && Y == 0) begin oled_data = 16'ha593; end
    else if (X == 10 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 11 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 12 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 13 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 14 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 15 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 16 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 17 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 18 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 19 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 20 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 21 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 22 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 23 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 24 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 25 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 26 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 27 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 28 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 29 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 30 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 31 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 32 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 33 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 34 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 35 && Y == 0) begin oled_data = 16'h84ce; end
    else if (X == 36 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 37 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 38 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 39 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 40 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 41 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 42 && Y == 0) begin oled_data = 16'h84ce; end
    else if (X == 43 && Y == 0) begin oled_data = 16'h84ce; end
    else if (X == 44 && Y == 0) begin oled_data = 16'h84ce; end
    else if (X == 45 && Y == 0) begin oled_data = 16'h84ce; end
    else if (X == 46 && Y == 0) begin oled_data = 16'h9cb1; end
    else if (X == 47 && Y == 0) begin oled_data = 16'hb573; end
    else if (X == 48 && Y == 0) begin oled_data = 16'hc5d4; end
    else if (X == 49 && Y == 0) begin oled_data = 16'had31; end
    else if (X == 50 && Y == 0) begin oled_data = 16'h84ce; end
    else if (X == 51 && Y == 0) begin oled_data = 16'h84ce; end
    else if (X == 52 && Y == 0) begin oled_data = 16'h84ce; end
    else if (X == 53 && Y == 0) begin oled_data = 16'h84ce; end
    else if (X == 54 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 55 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 56 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 57 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 58 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 59 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 60 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 61 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 62 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 63 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 64 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 65 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 66 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 67 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 68 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 69 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 70 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 71 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 72 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 73 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 74 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 75 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 76 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 77 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 78 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 79 && Y == 0) begin oled_data = 16'h84ce; end
    else if (X == 80 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 81 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 82 && Y == 0) begin oled_data = 16'h84ce; end
    else if (X == 83 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 84 && Y == 0) begin oled_data = 16'h84ce; end
    else if (X == 85 && Y == 0) begin oled_data = 16'had31; end
    else if (X == 86 && Y == 0) begin oled_data = 16'hc5d4; end
    else if (X == 87 && Y == 0) begin oled_data = 16'hb573; end
    else if (X == 88 && Y == 0) begin oled_data = 16'h84ce; end
    else if (X == 89 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 90 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 91 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 92 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 93 && Y == 0) begin oled_data = 16'h8d0f; end
    else if (X == 94 && Y == 0) begin oled_data = 16'h9551; end
    else if (X == 95 && Y == 0) begin oled_data = 16'hb5b6; end
    else if (X == 0 && Y == 1) begin oled_data = 16'h9551; end
    else if (X >= 1 && X <= 2 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 3 && Y == 1) begin oled_data = 16'h6468; end
    else if (X == 4 && Y == 1) begin oled_data = 16'h64a9; end
    else if (X == 5 && Y == 1) begin oled_data = 16'h6468; end
    else if (X == 6 && Y == 1) begin oled_data = 16'h6468; end
    else if (X == 7 && Y == 1) begin oled_data = 16'h6468; end
    else if (X == 8 && Y == 1) begin oled_data = 16'h6468; end
    else if (X == 9 && Y == 1) begin oled_data = 16'h6468; end
    else if (X == 10 && Y == 1) begin oled_data = 16'h6468; end
    else if (X == 11 && Y == 1) begin oled_data = 16'h6468; end
    else if (X == 12 && Y == 1) begin oled_data = 16'h6468; end
    else if (X >= 13 && X <= 15 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 16 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 17 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 18 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 19 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 20 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 21 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 22 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 23 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 24 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 25 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 26 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 27 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 28 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 29 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 30 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 31 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 32 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 33 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 34 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 35 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 36 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 37 && Y == 1) begin oled_data = 16'h4346; end
    else if (X == 38 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 39 && Y == 1) begin oled_data = 16'h4346; end
    else if (X == 40 && Y == 1) begin oled_data = 16'h4346; end
    else if (X == 41 && Y == 1) begin oled_data = 16'h4346; end
    else if (X == 42 && Y == 1) begin oled_data = 16'h4346; end
    else if (X == 43 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 44 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 45 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 46 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X == 47 && Y == 1) begin oled_data = 16'hcdd1; end
    else if (X == 49 && Y == 1) begin oled_data = 16'ha4ee; end
    else if (X == 50 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X >= 51 && X <= 52 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 53 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X >= 54 && X <= 59 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 60 && Y == 1) begin oled_data = 16'h6468; end
    else if (X == 61 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 62 && Y == 1) begin oled_data = 16'h6468; end
    else if (X >= 63 && X <= 64 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 65 && Y == 1) begin oled_data = 16'h6468; end
    else if (X >= 66 && X <= 68 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 69 && Y == 1) begin oled_data = 16'h53c7; end
    else if (X >= 70 && X <= 72 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 73 && Y == 1) begin oled_data = 16'h6468; end
    else if (X >= 74 && X <= 75 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 76 && Y == 1) begin oled_data = 16'h6468; end
    else if (X == 77 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 78 && Y == 1) begin oled_data = 16'h6468; end
    else if (X == 79 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 80 && Y == 1) begin oled_data = 16'h6468; end
    else if (X == 81 && Y == 1) begin oled_data = 16'h6468; end
    else if (X >= 82 && X <= 83 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 84 && Y == 1) begin oled_data = 16'h740a; end
    else if (X == 85 && Y == 1) begin oled_data = 16'hcdd1; end
    else if (X == 87 && Y == 1) begin oled_data = 16'ha4ee; end
    else if (X >= 88 && X <= 89 && Y == 1) begin oled_data = 16'h5c27; end
    else if (X == 90 && Y == 1) begin oled_data = 16'h6468; end
    else if (X == 91 && Y == 1) begin oled_data = 16'h6468; end
    else if (X == 92 && Y == 1) begin oled_data = 16'h64a9; end
    else if (X == 93 && Y == 1) begin oled_data = 16'h64a9; end
    else if (X == 94 && Y == 1) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 1) begin oled_data = 16'h8d0f; end
    else if (X == 0 && Y == 2) begin oled_data = 16'h9551; end
    else if (X == 1 && Y == 2) begin oled_data = 16'h6468; end
    else if (X == 2 && Y == 2) begin oled_data = 16'h5c27; end
    else if (X == 3 && Y == 2) begin oled_data = 16'h6468; end
    else if (X == 4 && Y == 2) begin oled_data = 16'h6468; end
    else if (X == 5 && Y == 2) begin oled_data = 16'h6468; end
    else if (X == 6 && Y == 2) begin oled_data = 16'h64a9; end
    else if (X == 7 && Y == 2) begin oled_data = 16'h64a9; end
    else if (X == 8 && Y == 2) begin oled_data = 16'h64a9; end
    else if (X == 9 && Y == 2) begin oled_data = 16'h64a9; end
    else if (X == 10 && Y == 2) begin oled_data = 16'h6468; end
    else if (X == 11 && Y == 2) begin oled_data = 16'h64a9; end
    else if (X == 12 && Y == 2) begin oled_data = 16'h6468; end
    else if (X == 13 && Y == 2) begin oled_data = 16'h53c7; end
    else if (X == 14 && Y == 2) begin oled_data = 16'h5c27; end
    else if (X == 15 && Y == 2) begin oled_data = 16'h4225; end
    else if (X == 16 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 17 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 18 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 19 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 20 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 21 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 22 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 23 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 24 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 25 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 26 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 27 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 28 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 29 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 30 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 31 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 32 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 33 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 34 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 35 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 36 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 37 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 38 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 39 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 40 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 41 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 42 && Y == 2) begin oled_data = 16'h4285; end
    else if (X == 43 && Y == 2) begin oled_data = 16'h4346; end
    else if (X == 44 && Y == 2) begin oled_data = 16'h53c7; end
    else if (X == 45 && Y == 2) begin oled_data = 16'h53c7; end
    else if (X == 46 && Y == 2) begin oled_data = 16'h53c7; end
    else if (X == 47 && Y == 2) begin oled_data = 16'h948d; end
    else if (X == 48 && Y == 2) begin oled_data = 16'hbd91; end
    else if (X == 49 && Y == 2) begin oled_data = 16'hcdd1; end
    else if (X == 50 && Y == 2) begin oled_data = 16'h5bc8; end
    else if (X == 51 && Y == 2) begin oled_data = 16'h53c7; end
    else if (X == 52 && Y == 2) begin oled_data = 16'h4346; end
    else if (X == 53 && Y == 2) begin oled_data = 16'h4225; end
    else if (X == 54 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 55 && Y == 2) begin oled_data = 16'h72e7; end
    else if (X == 56 && Y == 2) begin oled_data = 16'h72e7; end
    else if (X == 57 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 58 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 59 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 60 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 61 && Y == 2) begin oled_data = 16'h72e7; end
    else if (X == 62 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 63 && Y == 2) begin oled_data = 16'h72e7; end
    else if (X == 64 && Y == 2) begin oled_data = 16'h72e7; end
    else if (X == 65 && Y == 2) begin oled_data = 16'h72e7; end
    else if (X == 66 && Y == 2) begin oled_data = 16'h72e7; end
    else if (X == 67 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 68 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 69 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 70 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 71 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 72 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 73 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 74 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 75 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 76 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 77 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 78 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 79 && Y == 2) begin oled_data = 16'h6aa7; end
    else if (X == 80 && Y == 2) begin oled_data = 16'h53c7; end
    else if (X == 81 && Y == 2) begin oled_data = 16'h5c27; end
    else if (X == 82 && Y == 2) begin oled_data = 16'h53c7; end
    else if (X == 83 && Y == 2) begin oled_data = 16'h63e9; end
    else if (X >= 84 && X <= 86 && Y == 2) begin oled_data = 16'hcdd1; end
    else if (X == 87 && Y == 2) begin oled_data = 16'h5bc8; end
    else if (X >= 88 && X <= 89 && Y == 2) begin oled_data = 16'h5c27; end
    else if (X == 90 && Y == 2) begin oled_data = 16'h6468; end
    else if (X == 91 && Y == 2) begin oled_data = 16'h64a9; end
    else if (X == 92 && Y == 2) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 2) begin oled_data = 16'h64a9; end
    else if (X == 94 && Y == 2) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 2) begin oled_data = 16'h9551; end
    else if (X == 0 && Y == 3) begin oled_data = 16'h9551; end
    else if (X == 1 && Y == 3) begin oled_data = 16'h6468; end
    else if (X == 2 && Y == 3) begin oled_data = 16'h64a9; end
    else if (X == 3 && Y == 3) begin oled_data = 16'h64a9; end
    else if (X == 4 && Y == 3) begin oled_data = 16'h64a9; end
    else if (X == 5 && Y == 3) begin oled_data = 16'h7509; end
    else if (X == 6 && Y == 3) begin oled_data = 16'h7509; end
    else if (X == 7 && Y == 3) begin oled_data = 16'h64a9; end
    else if (X == 8 && Y == 3) begin oled_data = 16'h64a9; end
    else if (X == 9 && Y == 3) begin oled_data = 16'h64a9; end
    else if (X == 10 && Y == 3) begin oled_data = 16'h64a9; end
    else if (X == 11 && Y == 3) begin oled_data = 16'h64a9; end
    else if (X == 12 && Y == 3) begin oled_data = 16'h6468; end
    else if (X == 13 && Y == 3) begin oled_data = 16'h5c27; end
    else if (X == 14 && Y == 3) begin oled_data = 16'h53c7; end
    else if (X == 15 && Y == 3) begin oled_data = 16'h3263; end
    else if (X == 16 && Y == 3) begin oled_data = 16'h5a87; end
    else if (X == 17 && Y == 3) begin oled_data = 16'h6b4d; end
    else if (X == 18 && Y == 3) begin oled_data = 16'h6b4d; end
    else if (X >= 19 && X <= 38 && Y == 3) begin oled_data = 16'h8c71; end
    else if (X == 39 && Y == 3) begin oled_data = 16'h840f; end
    else if (X == 40 && Y == 3) begin oled_data = 16'h5b0c; end
    else if (X == 41 && Y == 3) begin oled_data = 16'h5b0c; end
    else if (X == 42 && Y == 3) begin oled_data = 16'h4225; end
    else if (X == 43 && Y == 3) begin oled_data = 16'h4346; end
    else if (X >= 44 && X <= 46 && Y == 3) begin oled_data = 16'h5c27; end
    else if (X == 47 && Y == 3) begin oled_data = 16'h53c7; end
    else if (X == 50 && Y == 3) begin oled_data = 16'h7c4b; end
    else if (X == 51 && Y == 3) begin oled_data = 16'h53c7; end
    else if (X == 52 && Y == 3) begin oled_data = 16'h4346; end
    else if (X == 53 && Y == 3) begin oled_data = 16'h39c5; end
    else if (X == 54 && Y == 3) begin oled_data = 16'h6b4d; end
    else if (X == 55 && Y == 3) begin oled_data = 16'h6b4d; end
    else if (X == 56 && Y == 3) begin oled_data = 16'h8c71; end
    else if (X == 57 && Y == 3) begin oled_data = 16'h94b2; end
    else if (X == 58 && Y == 3) begin oled_data = 16'h94b2; end
    else if (X == 59 && Y == 3) begin oled_data = 16'h94b2; end
    else if (X == 60 && Y == 3) begin oled_data = 16'h94b2; end
    else if (X == 61 && Y == 3) begin oled_data = 16'h94b2; end
    else if (X == 62 && Y == 3) begin oled_data = 16'h94b2; end
    else if (X == 63 && Y == 3) begin oled_data = 16'h94b2; end
    else if (X == 64 && Y == 3) begin oled_data = 16'h94b2; end
    else if (X == 65 && Y == 3) begin oled_data = 16'h94b2; end
    else if (X == 66 && Y == 3) begin oled_data = 16'h94b2; end
    else if (X == 67 && Y == 3) begin oled_data = 16'h8c71; end
    else if (X >= 68 && X <= 76 && Y == 3) begin oled_data = 16'h94b2; end
    else if (X == 77 && Y == 3) begin oled_data = 16'h6b4d; end
    else if (X == 78 && Y == 3) begin oled_data = 16'h6b4d; end
    else if (X == 79 && Y == 3) begin oled_data = 16'h4a27; end
    else if (X == 80 && Y == 3) begin oled_data = 16'h53c7; end
    else if (X == 81 && Y == 3) begin oled_data = 16'h5c27; end
    else if (X == 82 && Y == 3) begin oled_data = 16'h53c7; end
    else if (X == 83 && Y == 3) begin oled_data = 16'hb550; end
    else if (X == 85 && Y == 3) begin oled_data = 16'hbd91; end
    else if (X == 86 && Y == 3) begin oled_data = 16'h740a; end
    else if (X >= 87 && X <= 89 && Y == 3) begin oled_data = 16'h5c27; end
    else if (X == 90 && Y == 3) begin oled_data = 16'h64a9; end
    else if (X == 91 && Y == 3) begin oled_data = 16'h7509; end
    else if (X == 92 && Y == 3) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 3) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 3) begin oled_data = 16'h7509; end
    else if (X == 95 && Y == 3) begin oled_data = 16'h9551; end
    else if (X == 0 && Y == 4) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 4) begin oled_data = 16'h64a9; end
    else if (X == 2 && Y == 4) begin oled_data = 16'h5c27; end
    else if (X == 3 && Y == 4) begin oled_data = 16'h64a9; end
    else if (X == 4 && Y == 4) begin oled_data = 16'h6468; end
    else if (X == 5 && Y == 4) begin oled_data = 16'h64a9; end
    else if (X == 6 && Y == 4) begin oled_data = 16'h7509; end
    else if (X == 7 && Y == 4) begin oled_data = 16'h64a9; end
    else if (X == 8 && Y == 4) begin oled_data = 16'h6468; end
    else if (X == 9 && Y == 4) begin oled_data = 16'h6468; end
    else if (X == 10 && Y == 4) begin oled_data = 16'h5c27; end
    else if (X == 11 && Y == 4) begin oled_data = 16'h6468; end
    else if (X == 12 && Y == 4) begin oled_data = 16'h5c27; end
    else if (X == 13 && Y == 4) begin oled_data = 16'h53c7; end
    else if (X == 14 && Y == 4) begin oled_data = 16'h4346; end
    else if (X == 15 && Y == 4) begin oled_data = 16'h3263; end
    else if (X == 16 && Y == 4) begin oled_data = 16'h5a87; end
    else if (X == 17 && Y == 4) begin oled_data = 16'h6b4d; end
    else if (X == 18 && Y == 4) begin oled_data = 16'h73af; end
    else if (X >= 19 && X <= 38  && Y == 4) begin oled_data = 16'hbdd7; end
    else if (X == 39 && Y == 4) begin oled_data = 16'hb5b6; end
    else if (X == 40 && Y == 4) begin oled_data = 16'h6b4d; end
    else if (X == 41 && Y == 4) begin oled_data = 16'h5b0c; end
    else if (X == 42 && Y == 4) begin oled_data = 16'h4225; end
    else if (X == 43 && Y == 4) begin oled_data = 16'h4346; end
    else if (X == 44 && Y == 4) begin oled_data = 16'h53c7; end
    else if (X == 45 && Y == 4) begin oled_data = 16'h53c7; end
    else if (X == 46 && Y == 4) begin oled_data = 16'h53c7; end
    else if (X == 47 && Y == 4) begin oled_data = 16'h53c7; end
    else if (X == 48 && Y == 4) begin oled_data = 16'hcdd1; end
    else if (X == 50 && Y == 4) begin oled_data = 16'had0f; end
    else if (X == 51 && Y == 4) begin oled_data = 16'h5b88; end
    else if (X == 52 && Y == 4) begin oled_data = 16'h4346; end
    else if (X == 53 && Y == 4) begin oled_data = 16'h4225; end
    else if (X == 54 && Y == 4) begin oled_data = 16'h6b4d; end
    else if (X == 55 && Y == 4) begin oled_data = 16'h5b0c; end
    else if (X == 56 && Y == 4) begin oled_data = 16'had55; end
    else if (X == 57 && Y == 4) begin oled_data = 16'hb5b6; end
    else if (X == 58 && Y == 4) begin oled_data = 16'hb5b6; end
    else if (X == 59 && Y == 4) begin oled_data = 16'hb5b6; end
    else if (X == 60 && Y == 4) begin oled_data = 16'hbdd7; end
    else if (X == 61 && Y == 4) begin oled_data = 16'hbdd7; end
    else if (X == 62 && Y == 4) begin oled_data = 16'hb5b6; end
    else if (X == 63 && Y == 4) begin oled_data = 16'hb5b6; end
    else if (X == 64 && Y == 4) begin oled_data = 16'hb5b6; end
    else if (X == 65 && Y == 4) begin oled_data = 16'hbdd7; end
    else if (X == 66 && Y == 4) begin oled_data = 16'hbdd7; end
    else if (X == 67 && Y == 4) begin oled_data = 16'hbdd7; end
    else if (X == 68 && Y == 4) begin oled_data = 16'hb5b6; end
    else if (X == 69 && Y == 4) begin oled_data = 16'hb5b6; end
    else if (X == 70 && Y == 4) begin oled_data = 16'hb5b6; end
    else if (X == 71 && Y == 4) begin oled_data = 16'hbdd7; end
    else if (X == 72 && Y == 4) begin oled_data = 16'hb5b6; end
    else if (X == 73 && Y == 4) begin oled_data = 16'hb5b6; end
    else if (X == 74 && Y == 4) begin oled_data = 16'hbdd7; end
    else if (X == 75 && Y == 4) begin oled_data = 16'hbdd7; end
    else if (X == 76 && Y == 4) begin oled_data = 16'hb5b6; end
    else if (X == 77 && Y == 4) begin oled_data = 16'h73af; end
    else if (X == 78 && Y == 4) begin oled_data = 16'h6b4d; end
    else if (X == 79 && Y == 4) begin oled_data = 16'h4a27; end
    else if (X == 80 && Y == 4) begin oled_data = 16'h53c7; end
    else if (X == 81 && Y == 4) begin oled_data = 16'h5c27; end
    else if (X == 82 && Y == 4) begin oled_data = 16'h5bc8; end
    else if (X == 83 && Y == 4) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 4) begin oled_data = 16'ha4ee; end
    else if (X == 86 && Y == 4) begin oled_data = 16'h53c7; end
    else if (X == 87 && Y == 4) begin oled_data = 16'h53c7; end
    else if (X >= 88 && X <= 89 && Y == 4) begin oled_data = 16'h5c27; end
    else if (X == 90 && Y == 4) begin oled_data = 16'h6468; end
    else if (X == 91 && Y == 4) begin oled_data = 16'h7509; end
    else if (X == 92 && Y == 4) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 4) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 4) begin oled_data = 16'h7509; end
    else if (X == 95 && Y == 4) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 5) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 5) begin oled_data = 16'h6468; end
    else if (X == 2 && Y == 5) begin oled_data = 16'h64a9; end
    else if (X == 3 && Y == 5) begin oled_data = 16'h6468; end
    else if (X == 4 && Y == 5) begin oled_data = 16'h6468; end
    else if (X == 5 && Y == 5) begin oled_data = 16'h6468; end
    else if (X == 6 && Y == 5) begin oled_data = 16'h64a9; end
    else if (X == 7 && Y == 5) begin oled_data = 16'h64a9; end
    else if (X == 8 && Y == 5) begin oled_data = 16'h64a9; end
    else if (X == 9 && Y == 5) begin oled_data = 16'h6468; end
    else if (X >= 10 && X <= 12 && Y == 5) begin oled_data = 16'h5c27; end
    else if (X == 13 && Y == 5) begin oled_data = 16'h4346; end
    else if (X == 14 && Y == 5) begin oled_data = 16'h4346; end
    else if (X == 15 && Y == 5) begin oled_data = 16'h3263; end
    else if (X == 16 && Y == 5) begin oled_data = 16'h5a87; end
    else if (X == 17 && Y == 5) begin oled_data = 16'h6b4d; end
    else if (X == 18 && Y == 5) begin oled_data = 16'h73af; end
    else if (X == 19 && Y == 5) begin oled_data = 16'ha514; end
    else if (X >= 20 && X <= 38  && Y == 5) begin oled_data = 16'ha514; end
    else if (X == 39 && Y == 5) begin oled_data = 16'h94b2; end
    else if (X == 40 && Y == 5) begin oled_data = 16'h5b0c; end
    else if (X == 41 && Y == 5) begin oled_data = 16'h5b0c; end
    else if (X == 42 && Y == 5) begin oled_data = 16'h4225; end
    else if (X == 43 && Y == 5) begin oled_data = 16'h848c; end
    else if (X >= 44 && X <= 50 && Y == 5) begin oled_data = 16'hcdd1; end
    else if (X == 52 && Y == 5) begin oled_data = 16'h948d; end
    else if (X == 53 && Y == 5) begin oled_data = 16'h39c5; end
    else if (X == 54 && Y == 5) begin oled_data = 16'h5b0c; end
    else if (X == 55 && Y == 5) begin oled_data = 16'h5b0c; end
    else if (X == 56 && Y == 5) begin oled_data = 16'h94b2; end
    else if (X >= 57 && X <= 71 && Y == 5) begin oled_data = 16'ha514; end
    else if (X == 72 && Y == 5) begin oled_data = 16'had55; end
    else if (X == 73 && Y == 5) begin oled_data = 16'ha514; end
    else if (X == 74 && Y == 5) begin oled_data = 16'ha514; end
    else if (X == 75 && Y == 5) begin oled_data = 16'ha514; end
    else if (X == 76 && Y == 5) begin oled_data = 16'ha514; end
    else if (X == 77 && Y == 5) begin oled_data = 16'h6b4d; end
    else if (X == 78 && Y == 5) begin oled_data = 16'h5b0c; end
    else if (X == 79 && Y == 5) begin oled_data = 16'h4a27; end
    else if (X == 80 && Y == 5) begin oled_data = 16'h53c7; end
    else if (X == 81 && Y == 5) begin oled_data = 16'h5c27; end
    else if (X == 82 && Y == 5) begin oled_data = 16'h740a; end
    else if (X == 85 && Y == 5) begin oled_data = 16'h948d; end
    else if (X >= 86 && X <= 89 && Y == 5) begin oled_data = 16'h5c27; end
    else if (X == 90 && Y == 5) begin oled_data = 16'h6468; end
    else if (X == 91 && Y == 5) begin oled_data = 16'h7509; end
    else if (X == 92 && Y == 5) begin oled_data = 16'h7d6b; end
    else if (X == 93 && Y == 5) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 5) begin oled_data = 16'h7509; end
    else if (X == 95 && Y == 5) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 6) begin oled_data = 16'ha593; end
    else if (X >= 1 && X <= 8 && Y == 6) begin oled_data = 16'h5c27; end
    else if (X == 9 && Y == 6) begin oled_data = 16'h6468; end
    else if (X >= 10 && X <= 11 && Y == 6) begin oled_data = 16'h5c27; end
    else if (X == 12 && Y == 6) begin oled_data = 16'h53c7; end
    else if (X == 13 && Y == 6) begin oled_data = 16'h4346; end
    else if (X == 14 && Y == 6) begin oled_data = 16'h4346; end
    else if (X == 15 && Y == 6) begin oled_data = 16'h3263; end
    else if (X == 16 && Y == 6) begin oled_data = 16'h5a87; end
    else if (X == 17 && Y == 6) begin oled_data = 16'h5b0c; end
    else if (X == 18 && Y == 6) begin oled_data = 16'h73af; end
    else if (X == 19 && Y == 6) begin oled_data = 16'hb5b6; end
    else if (X == 20 && Y == 6) begin oled_data = 16'hbdd7; end
    else if (X == 21 && Y == 6) begin oled_data = 16'hbdd7; end
    else if (X >= 22 && X <= 38 && Y == 6) begin oled_data = 16'hb5b6; end
    else if (X == 39 && Y == 6) begin oled_data = 16'had55; end
    else if (X == 40 && Y == 6) begin oled_data = 16'h5b0c; end
    else if (X == 41 && Y == 6) begin oled_data = 16'h52ca; end
    else if (X == 42 && Y == 6) begin oled_data = 16'h5a87; end
    else if (X == 50 && Y == 6) begin oled_data = 16'hcdd1; end
    else if (X == 52 && Y == 6) begin oled_data = 16'had0f; end
    else if (X == 53 && Y == 6) begin oled_data = 16'h39c5; end
    else if (X == 54 && Y == 6) begin oled_data = 16'h52ca; end
    else if (X == 55 && Y == 6) begin oled_data = 16'h52ca; end
    else if (X == 56 && Y == 6) begin oled_data = 16'had55; end
    else if (X == 57 && Y == 6) begin oled_data = 16'hb5b6; end
    else if (X == 58 && Y == 6) begin oled_data = 16'hbdd7; end
    else if (X >= 59 && X <= 71 &&  Y == 6) begin oled_data = 16'hb5b6; end
    else if (X == 72 && Y == 6) begin oled_data = 16'hbdd7; end
    else if (X == 73 && Y == 6) begin oled_data = 16'hbdd7; end
    else if (X == 74 && Y == 6) begin oled_data = 16'hbdd7; end
    else if (X == 75 && Y == 6) begin oled_data = 16'hb5b6; end
    else if (X == 76 && Y == 6) begin oled_data = 16'hb5b6; end
    else if (X == 77 && Y == 6) begin oled_data = 16'h6b4d; end
    else if (X == 78 && Y == 6) begin oled_data = 16'h5b0c; end
    else if (X == 79 && Y == 6) begin oled_data = 16'h4225; end
    else if (X == 80 && Y == 6) begin oled_data = 16'h4346; end
    else if (X == 81 && Y == 6) begin oled_data = 16'h53c7; end
    else if (X == 82 && Y == 6) begin oled_data = 16'h9cad; end
    else if (X == 85 && Y == 6) begin oled_data = 16'h740a; end
    else if (X >= 86 && X <= 88 && Y == 6) begin oled_data = 16'h5c27; end
    else if (X == 89 && Y == 6) begin oled_data = 16'h64a9; end
    else if (X == 90 && Y == 6) begin oled_data = 16'h7509; end
    else if (X == 91 && Y == 6) begin oled_data = 16'h7509; end
    else if (X == 92 && Y == 6) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 6) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 6) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 6) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 7) begin oled_data = 16'h9551; end
    else if (X == 1 && Y == 7) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 7) begin oled_data = 16'h4b07; end
    else if (X == 3 && Y == 7) begin oled_data = 16'h4285; end
    else if (X == 4 && Y == 7) begin oled_data = 16'h4285; end
    else if (X == 5 && Y == 7) begin oled_data = 16'h4225; end
    else if (X == 6 && Y == 7) begin oled_data = 16'h4225; end
    else if (X == 7 && Y == 7) begin oled_data = 16'h4225; end
    else if (X == 8 && Y == 7) begin oled_data = 16'h4225; end
    else if (X == 9 && Y == 7) begin oled_data = 16'h4285; end
    else if (X == 10 && Y == 7) begin oled_data = 16'h4285; end
    else if (X == 11 && Y == 7) begin oled_data = 16'h53c7; end
    else if (X == 12 && Y == 7) begin oled_data = 16'h53c7; end
    else if (X == 13 && Y == 7) begin oled_data = 16'h4346; end
    else if (X == 14 && Y == 7) begin oled_data = 16'h63e9; end
    else if (X == 15 && Y == 7) begin oled_data = 16'h62e8; end
    else if (X == 16 && Y == 7) begin oled_data = 16'h4a27; end
    else if (X == 17 && Y == 7) begin oled_data = 16'h5b0c; end
    else if (X == 18 && Y == 7) begin oled_data = 16'h5b0c; end
    else if (X >= 19 && X <= 37 && Y == 7) begin oled_data = 16'h8c71; end
    else if (X == 38 && Y == 7) begin oled_data = 16'h94b2; end
    else if (X == 39 && Y == 7) begin oled_data = 16'h840f; end
    else if (X == 40 && Y == 7) begin oled_data = 16'h52ca; end
    else if (X == 41 && Y == 7) begin oled_data = 16'h4a89; end
    else if (X == 42 && Y == 7) begin oled_data = 16'h5a87; end
    else if (X >= 43 && X <= 44 && Y == 7) begin oled_data = 16'hcdd1; end
    else if (X == 45 && Y == 7) begin oled_data = 16'h840d; end
    else if (X == 46 && Y == 7) begin oled_data = 16'hb550; end
    else if (X == 47 && Y == 7) begin oled_data = 16'hb550; end
    else if (X == 48 && Y == 7) begin oled_data = 16'hb550; end
    else if (X == 49 && Y == 7) begin oled_data = 16'hb550; end
    else if (X == 50 && Y == 7) begin oled_data = 16'h840d; end
    else if (X == 51 && Y == 7) begin oled_data = 16'hcdd1; end
    else if (X == 52 && Y == 7) begin oled_data = 16'had0f; end
    else if (X == 53 && Y == 7) begin oled_data = 16'h39c5; end
    else if (X == 54 && Y == 7) begin oled_data = 16'h52ca; end
    else if (X == 55 && Y == 7) begin oled_data = 16'h4a89; end
    else if (X == 56 && Y == 7) begin oled_data = 16'h840f; end
    else if (X == 57 && Y == 7) begin oled_data = 16'h8c71; end
    else if (X == 58 && Y == 7) begin oled_data = 16'h94b2; end
    else if (X == 59 && Y == 7) begin oled_data = 16'h8c71; end
    else if (X == 60 && Y == 7) begin oled_data = 16'h8c71; end
    else if (X == 61 && Y == 7) begin oled_data = 16'h8c71; end
    else if (X == 62 && Y == 7) begin oled_data = 16'h8c71; end
    else if (X == 63 && Y == 7) begin oled_data = 16'h8c71; end
    else if (X == 64 && Y == 7) begin oled_data = 16'h8c71; end
    else if (X == 65 && Y == 7) begin oled_data = 16'h8c71; end
    else if (X == 66 && Y == 7) begin oled_data = 16'h8c71; end
    else if (X == 67 && Y == 7) begin oled_data = 16'h8c71; end
    else if (X == 68 && Y == 7) begin oled_data = 16'h8c71; end
    else if (X == 69 && Y == 7) begin oled_data = 16'h94b2; end
    else if (X == 70 && Y == 7) begin oled_data = 16'h8c71; end
    else if (X == 71 && Y == 7) begin oled_data = 16'h94b2; end
    else if (X == 72 && Y == 7) begin oled_data = 16'h94b2; end
    else if (X == 73 && Y == 7) begin oled_data = 16'ha514; end
    else if (X == 74 && Y == 7) begin oled_data = 16'h94b2; end
    else if (X == 75 && Y == 7) begin oled_data = 16'h94b2; end
    else if (X == 76 && Y == 7) begin oled_data = 16'h8c71; end
    else if (X == 77 && Y == 7) begin oled_data = 16'h5b0c; end
    else if (X == 78 && Y == 7) begin oled_data = 16'h5b0c; end
    else if (X == 79 && Y == 7) begin oled_data = 16'h4225; end
    else if (X == 80 && Y == 7) begin oled_data = 16'h7c4b; end
    else if (X == 81 && Y == 7) begin oled_data = 16'had0f; end
    else if (X == 82 && Y == 7) begin oled_data = 16'hbd91; end
    else if (X == 85 && Y == 7) begin oled_data = 16'had0f; end
    else if (X == 86 && Y == 7) begin oled_data = 16'h63e9; end
    else if (X == 87 && Y == 7) begin oled_data = 16'h5c27; end
    else if (X == 88 && Y == 7) begin oled_data = 16'h6468; end
    else if (X == 89 && Y == 7) begin oled_data = 16'h64a9; end
    else if (X == 90 && Y == 7) begin oled_data = 16'h64a9; end
    else if (X == 91 && Y == 7) begin oled_data = 16'h7509; end
    else if (X == 92 && Y == 7) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 7) begin oled_data = 16'h64a9; end
    else if (X == 94 && Y == 7) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 7) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 8) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 8) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 8) begin oled_data = 16'h4b07; end
    else if (X == 3 && Y == 8) begin oled_data = 16'h52ca; end
    else if (X == 4 && Y == 8) begin oled_data = 16'h840f; end
    else if (X == 5 && Y == 8) begin oled_data = 16'h4b0a; end
    else if (X == 6 && Y == 8) begin oled_data = 16'h4a89; end
    else if (X == 7 && Y == 8) begin oled_data = 16'h4b0a; end
    else if (X == 8 && Y == 8) begin oled_data = 16'h4b0a; end
    else if (X == 9 && Y == 8) begin oled_data = 16'h5a87; end
    else if (X == 10 && Y == 8) begin oled_data = 16'h4225; end
    else if (X == 11 && Y == 8) begin oled_data = 16'h5c27; end
    else if (X == 12 && Y == 8) begin oled_data = 16'h53c7; end
    else if (X == 13 && Y == 8) begin oled_data = 16'h9cad; end
    else if (X == 14 && Y == 8) begin oled_data = 16'hcd8f; end
    else if (X == 15 && Y == 8) begin oled_data = 16'h940c; end
    else if (X == 16 && Y == 8) begin oled_data = 16'h4a27; end
    else if (X == 17 && Y == 8) begin oled_data = 16'h52ca; end
    else if (X == 18 && Y == 8) begin oled_data = 16'h5b0c; end
    else if (X >= 19 && X <= 33 && Y == 8) begin oled_data = 16'ha514; end
    else if (X == 34 && Y == 8) begin oled_data = 16'had55; end
    else if (X == 35 && Y == 8) begin oled_data = 16'had55; end
    else if (X == 36 && Y == 8) begin oled_data = 16'had55; end
    else if (X == 37 && Y == 8) begin oled_data = 16'had55; end
    else if (X == 38 && Y == 8) begin oled_data = 16'had55; end
    else if (X == 39 && Y == 8) begin oled_data = 16'h94b2; end
    else if (X == 40 && Y == 8) begin oled_data = 16'h4a89; end
    else if (X == 41 && Y == 8) begin oled_data = 16'h4a89; end
    else if (X == 42 && Y == 8) begin oled_data = 16'h5a87; end
    else if (X == 45 && Y == 8) begin oled_data = 16'hb550; end
    else if (X == 50 && Y == 8) begin oled_data = 16'had0f; end
    else if (X == 51 && Y == 8) begin oled_data = 16'hcdd1; end
    else if (X == 52 && Y == 8) begin oled_data = 16'had0f; end
    else if (X == 53 && Y == 8) begin oled_data = 16'h39c5; end
    else if (X == 54 && Y == 8) begin oled_data = 16'h4a89; end
    else if (X == 55 && Y == 8) begin oled_data = 16'h4a89; end
    else if (X == 56 && Y == 8) begin oled_data = 16'ha514; end
    else if (X >= 57 && X <= 76 && Y == 8) begin oled_data = 16'had55; end
    else if (X == 77 && Y == 8) begin oled_data = 16'h5b0c; end
    else if (X == 78 && Y == 8) begin oled_data = 16'h4a89; end
    else if (X == 79 && Y == 8) begin oled_data = 16'h39c5; end
    else if (X == 80 && Y == 8) begin oled_data = 16'had0f; end
    else if (X == 86 && Y == 8) begin oled_data = 16'hbd91; end
    else if (X == 87 && Y == 8) begin oled_data = 16'h53c7; end
    else if (X == 88 && Y == 8) begin oled_data = 16'h6468; end
    else if (X == 89 && Y == 8) begin oled_data = 16'h7509; end
    else if (X == 90 && Y == 8) begin oled_data = 16'h7509; end
    else if (X == 91 && Y == 8) begin oled_data = 16'h7509; end
    else if (X == 92 && Y == 8) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 8) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 8) begin oled_data = 16'h7509; end
    else if (X == 95 && Y == 8) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 9) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 9) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 9) begin oled_data = 16'h4b07; end
    else if (X == 3 && Y == 9) begin oled_data = 16'h52ca; end
    else if (X == 4 && Y == 9) begin oled_data = 16'h5bcd; end
    else if (X == 5 && Y == 9) begin oled_data = 16'h4b0a; end
    else if (X == 6 && Y == 9) begin oled_data = 16'h4b0a; end
    else if (X == 7 && Y == 9) begin oled_data = 16'h538c; end
    else if (X == 8 && Y == 9) begin oled_data = 16'h538c; end
    else if (X == 9 && Y == 9) begin oled_data = 16'h6b4a; end
    else if (X == 10 && Y == 9) begin oled_data = 16'h4285; end
    else if (X == 11 && Y == 9) begin oled_data = 16'h740a; end
    else if (X == 12 && Y == 9) begin oled_data = 16'h848c; end
    else if (X == 13 && Y == 9) begin oled_data = 16'had0f; end
    else if (X == 14 && Y == 9) begin oled_data = 16'hcd8f; end
    else if (X == 15 && Y == 9) begin oled_data = 16'h940c; end
    else if (X == 16 && Y == 9) begin oled_data = 16'h5a87; end
    else if (X == 17 && Y == 9) begin oled_data = 16'h940c; end
    else if (X == 18 && Y == 9) begin oled_data = 16'h83cc; end
    else if (X >= 19 && X <= 39 && Y == 9) begin oled_data = 16'h8c71; end
    else if (X == 40 && Y == 9) begin oled_data = 16'h83cc; end
    else if (X == 41 && Y == 9) begin oled_data = 16'h83cc; end
    else if (X == 42 && Y == 9) begin oled_data = 16'h5a87; end
    else if (X >= 43 && X <= 44 && Y == 9) begin oled_data = 16'hcdd1; end
    else if (X == 45 && Y == 9) begin oled_data = 16'had0f; end
    else if (X == 47 && Y == 9) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 9) begin oled_data = 16'hbd91; end
    else if (X == 49 && Y == 9) begin oled_data = 16'hcdd1; end
    else if (X == 50 && Y == 9) begin oled_data = 16'h9c8e; end
    else if (X == 51 && Y == 9) begin oled_data = 16'hcd8f; end
    else if (X == 52 && Y == 9) begin oled_data = 16'had0f; end
    else if (X == 53 && Y == 9) begin oled_data = 16'h39c5; end
    else if (X == 54 && Y == 9) begin oled_data = 16'h83cc; end
    else if (X == 55 && Y == 9) begin oled_data = 16'h83cc; end
    else if (X >= 56 && X <= 76&& Y == 9) begin oled_data = 16'h8c71; end
    else if (X == 77 && Y == 9) begin oled_data = 16'h83cc; end
    else if (X == 78 && Y == 9) begin oled_data = 16'h940c; end
    else if (X == 79 && Y == 9) begin oled_data = 16'h4225; end
    else if (X == 80 && Y == 9) begin oled_data = 16'hbd91; end
    else if (X == 82 && Y == 9) begin oled_data = 16'ha4f0; end
    else if (X == 83 && Y == 9) begin oled_data = 16'hb550; end
    else if (X == 84 && Y == 9) begin oled_data = 16'hb550; end
    else if (X == 85 && Y == 9) begin oled_data = 16'ha4f0; end
    else if (X == 86 && Y == 9) begin oled_data = 16'hcdd1; end
    else if (X == 87 && Y == 9) begin oled_data = 16'ha4ee; end
    else if (X == 88 && Y == 9) begin oled_data = 16'h5c27; end
    else if (X == 89 && Y == 9) begin oled_data = 16'h6468; end
    else if (X == 90 && Y == 9) begin oled_data = 16'h64a9; end
    else if (X == 91 && Y == 9) begin oled_data = 16'h64a9; end
    else if (X == 92 && Y == 9) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 9) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 9) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 9) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 10) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 10) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 10) begin oled_data = 16'h4285; end
    else if (X == 3 && Y == 10) begin oled_data = 16'h52ca; end
    else if (X == 4 && Y == 10) begin oled_data = 16'h5bcd; end
    else if (X == 5 && Y == 10) begin oled_data = 16'h4b0a; end
    else if (X == 6 && Y == 10) begin oled_data = 16'h4b0a; end
    else if (X == 7 && Y == 10) begin oled_data = 16'h5bcd; end
    else if (X == 8 && Y == 10) begin oled_data = 16'h5bcd; end
    else if (X == 9 && Y == 10) begin oled_data = 16'h6b4a; end
    else if (X == 10 && Y == 10) begin oled_data = 16'h62e8; end
    else if (X >= 13 && X <= 14 && Y == 10) begin oled_data = 16'hcdd1; end
    else if (X == 15 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 16 && Y == 10) begin oled_data = 16'hb550; end
    else if (X == 17 && Y == 10) begin oled_data = 16'hcdd1; end
    else if (X == 18 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 19 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 20 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 21 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 22 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 23 && Y == 10) begin oled_data = 16'hcdd1; end
    else if (X == 24 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 25 && Y == 10) begin oled_data = 16'hcdd1; end
    else if (X == 26 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 27 && Y == 10) begin oled_data = 16'hcdd1; end
    else if (X == 28 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 29 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 30 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 31 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 32 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 33 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 34 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X >= 35 && X <= 38 && Y == 10) begin oled_data = 16'hcdd1; end
    else if (X == 39 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 40 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 41 && Y == 10) begin oled_data = 16'hcdd1; end
    else if (X == 42 && Y == 10) begin oled_data = 16'hbd91; end
    else if (X == 45 && Y == 10) begin oled_data = 16'hb550; end
    else if (X == 47 && Y == 10) begin oled_data = 16'hbd91; end
    else if (X == 48 && Y == 10) begin oled_data = 16'hcdd1; end
    else if (X == 50 && Y == 10) begin oled_data = 16'hbd91; end
    else if (X >= 51 && X <= 52 && Y == 10) begin oled_data = 16'hcdd1; end
    else if (X == 53 && Y == 10) begin oled_data = 16'hb550; end
    else if (X == 54 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 55 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 56 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 57 && Y == 10) begin oled_data = 16'hcdd1; end
    else if (X == 58 && Y == 10) begin oled_data = 16'hb550; end
    else if (X == 59 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X == 60 && Y == 10) begin oled_data = 16'hcdd1; end
    else if (X >= 61 && X <= 77 && Y == 10) begin oled_data = 16'hcd8f; end
    else if (X >= 78 && X <= 82 && Y == 10) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 10) begin oled_data = 16'ha4f0; end
    else if (X == 88 && Y == 10) begin oled_data = 16'h5c27; end
    else if (X == 89 && Y == 10) begin oled_data = 16'h6468; end
    else if (X == 90 && Y == 10) begin oled_data = 16'h64a9; end
    else if (X == 91 && Y == 10) begin oled_data = 16'h7509; end
    else if (X == 92 && Y == 10) begin oled_data = 16'h7d6b; end
    else if (X == 93 && Y == 10) begin oled_data = 16'h7d6b; end
    else if (X == 94 && Y == 10) begin oled_data = 16'h7d6b; end
    else if (X == 95 && Y == 10) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 11) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 11) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 11) begin oled_data = 16'h4b07; end
    else if (X == 3 && Y == 11) begin oled_data = 16'h52ca; end
    else if (X == 4 && Y == 11) begin oled_data = 16'h840f; end
    else if (X == 5 && Y == 11) begin oled_data = 16'h4b0a; end
    else if (X == 6 && Y == 11) begin oled_data = 16'h4b0a; end
    else if (X == 7 && Y == 11) begin oled_data = 16'h5bcd; end
    else if (X == 8 && Y == 11) begin oled_data = 16'h538c; end
    else if (X == 9 && Y == 11) begin oled_data = 16'h62e8; end
    else if (X == 10 && Y == 11) begin oled_data = 16'h62e8; end
    else if (X >= 13 && X <= 25 && Y == 11) begin oled_data = 16'hcdd1; end
    else if (X == 26 && Y == 11) begin oled_data = 16'hcd8f; end
    else if (X >= 27 && X <= 42 && Y == 11) begin oled_data = 16'hcdd1; end
    else if (X == 45 && Y == 11) begin oled_data = 16'had0f; end
    else if (X >= 47 && X <= 57 && Y == 11) begin oled_data = 16'hcdd1; end
    else if (X == 58 && Y == 11) begin oled_data = 16'hcd8f; end
    else if (X >= 59 && X <= 62 && Y == 11) begin oled_data = 16'hcdd1; end
    else if (X == 63 && Y == 11) begin oled_data = 16'hcd8f; end
    else if (X >= 64 && X <= 79 && Y == 11) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 11) begin oled_data = 16'hb550; end
    else if (X == 88 && Y == 11) begin oled_data = 16'h740a; end
    else if (X == 89 && Y == 11) begin oled_data = 16'h6468; end
    else if (X == 90 && Y == 11) begin oled_data = 16'h64a9; end
    else if (X == 91 && Y == 11) begin oled_data = 16'h7509; end
    else if (X == 92 && Y == 11) begin oled_data = 16'h7d6b; end
    else if (X == 93 && Y == 11) begin oled_data = 16'h7d6b; end
    else if (X == 94 && Y == 11) begin oled_data = 16'h7d6b; end
    else if (X == 95 && Y == 11) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 12) begin oled_data = 16'h9551; end
    else if (X == 1 && Y == 12) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 12) begin oled_data = 16'h4285; end
    else if (X == 3 && Y == 12) begin oled_data = 16'h4a89; end
    else if (X == 4 && Y == 12) begin oled_data = 16'h538c; end
    else if (X == 5 && Y == 12) begin oled_data = 16'h4b0a; end
    else if (X == 6 && Y == 12) begin oled_data = 16'h4b0a; end
    else if (X == 7 && Y == 12) begin oled_data = 16'h538c; end
    else if (X == 8 && Y == 12) begin oled_data = 16'h538c; end
    else if (X == 9 && Y == 12) begin oled_data = 16'h538c; end
    else if (X == 10 && Y == 12) begin oled_data = 16'h62e8; end
    else if (X >= 11 && X <= 12 && Y == 12) begin oled_data = 16'hcdd1; end
    else if (X == 13 && Y == 12) begin oled_data = 16'h83cc; end
    else if (X >= 14 && X <= 26 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 27 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 28 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 29 && Y == 12) begin oled_data = 16'h948d; end
    else if (X == 30 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 31 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 32 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 33 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 34 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 35 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 36 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 37 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 38 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 39 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 40 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 41 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 42 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 43 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 44 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 45 && Y == 12) begin oled_data = 16'h9c8e; end
    else if (X == 47 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 48 && Y == 12) begin oled_data = 16'ha4f0; end
    else if (X == 49 && Y == 12) begin oled_data = 16'hbd91; end
    else if (X == 50 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 51 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 52 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 53 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 54 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 55 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 56 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 57 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 58 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 59 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 60 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 61 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 62 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 63 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 64 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 65 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 66 && Y == 12) begin oled_data = 16'h9c8e; end
    else if (X == 67 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 68 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 69 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 70 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 71 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 72 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 73 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 74 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 75 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 76 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 77 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 78 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 79 && Y == 12) begin oled_data = 16'had0f; end
    else if (X == 80 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 81 && Y == 12) begin oled_data = 16'hb550; end
    else if (X == 82 && Y == 12) begin oled_data = 16'h9c8e; end
    else if (X == 85 && Y == 12) begin oled_data = 16'ha4f0; end
    else if (X == 87 && Y == 12) begin oled_data = 16'hcdd1; end
    else if (X == 88 && Y == 12) begin oled_data = 16'h740a; end
    else if (X == 89 && Y == 12) begin oled_data = 16'h5c27; end
    else if (X == 90 && Y == 12) begin oled_data = 16'h64a9; end
    else if (X == 91 && Y == 12) begin oled_data = 16'h7d6b; end
    else if (X == 92 && Y == 12) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 12) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 12) begin oled_data = 16'h7509; end
    else if (X == 95 && Y == 12) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 13) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 13) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 13) begin oled_data = 16'h4285; end
    else if (X == 3 && Y == 13) begin oled_data = 16'h5b0c; end
    else if (X == 4 && Y == 13) begin oled_data = 16'h8c71; end
    else if (X == 5 && Y == 13) begin oled_data = 16'h4b0a; end
    else if (X == 6 && Y == 13) begin oled_data = 16'h4b0a; end
    else if (X == 7 && Y == 13) begin oled_data = 16'h5bcd; end
    else if (X == 8 && Y == 13) begin oled_data = 16'h5bcd; end
    else if (X == 9 && Y == 13) begin oled_data = 16'h538c; end
    else if (X == 10 && Y == 13) begin oled_data = 16'h6b4a; end
    else if (X == 13 && Y == 13) begin oled_data = 16'had0f; end
    else if (X >= 26 && X <= 56 && Y == 13) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 13) begin oled_data = 16'hb550; end
    else if (X == 88 && Y == 13) begin oled_data = 16'h7c4b; end
    else if (X == 89 && Y == 13) begin oled_data = 16'h5c27; end
    else if (X == 90 && Y == 13) begin oled_data = 16'h64a9; end
    else if (X == 91 && Y == 13) begin oled_data = 16'h7509; end
    else if (X == 92 && Y == 13) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 13) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 13) begin oled_data = 16'h7509; end
    else if (X == 95 && Y == 13) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 14) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 14) begin oled_data = 16'h53c7; end
    else if (X == 2 && Y == 14) begin oled_data = 16'h4285; end
    else if (X == 3 && Y == 14) begin oled_data = 16'h39c5; end
    else if (X == 4 && Y == 14) begin oled_data = 16'h39c5; end
    else if (X == 5 && Y == 14) begin oled_data = 16'h39c5; end
    else if (X == 6 && Y == 14) begin oled_data = 16'h39c5; end
    else if (X == 7 && Y == 14) begin oled_data = 16'h39c5; end
    else if (X == 8 && Y == 14) begin oled_data = 16'h39c5; end
    else if (X == 9 && Y == 14) begin oled_data = 16'h39c5; end
    else if (X == 10 && Y == 14) begin oled_data = 16'h5a87; end
    else if (X == 11 && Y == 14) begin oled_data = 16'hcdd1; end
    else if (X == 13 && Y == 14) begin oled_data = 16'had0f; end
    else if (X == 15 && Y == 14) begin oled_data = 16'hbd91; end
    else if (X == 16 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 17 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 18 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 19 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 20 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 21 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 22 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 23 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 24 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 25 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 26 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 27 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 28 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 29 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 30 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 31 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 32 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 33 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 34 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 35 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 36 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 37 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 38 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 39 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 40 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 41 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 42 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 43 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 44 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 45 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 46 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 47 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 48 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 49 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 50 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 51 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 52 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 53 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 54 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 55 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 56 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 57 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 58 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 59 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 60 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 61 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 62 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 63 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 64 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 65 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 66 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 67 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 68 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 69 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 70 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 71 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 72 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 73 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 74 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 75 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 76 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 77 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 78 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 79 && Y == 14) begin oled_data = 16'had31; end
    else if (X == 80 && Y == 14) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 14) begin oled_data = 16'ha4f0; end
    else if (X == 83 && Y == 14) begin oled_data = 16'hb550; end
    else if (X == 84 && Y == 14) begin oled_data = 16'hb550; end
    else if (X == 85 && Y == 14) begin oled_data = 16'h9c8e; end
    else if (X == 87 && Y == 14) begin oled_data = 16'hcdd1; end
    else if (X == 88 && Y == 14) begin oled_data = 16'h63e9; end
    else if (X >= 89 && X <= 90 && Y == 14) begin oled_data = 16'h5c27; end
    else if (X == 91 && Y == 14) begin oled_data = 16'h64a9; end
    else if (X == 92 && Y == 14) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 14) begin oled_data = 16'h64a9; end
    else if (X == 94 && Y == 14) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 14) begin oled_data = 16'h9551; end
    else if (X == 0 && Y == 15) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 15) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 15) begin oled_data = 16'h4285; end
    else if (X == 3 && Y == 15) begin oled_data = 16'h4a89; end
    else if (X == 4 && Y == 15) begin oled_data = 16'h538c; end
    else if (X == 5 && Y == 15) begin oled_data = 16'h4b0a; end
    else if (X == 6 && Y == 15) begin oled_data = 16'h4b0a; end
    else if (X == 7 && Y == 15) begin oled_data = 16'h538c; end
    else if (X == 8 && Y == 15) begin oled_data = 16'h538c; end
    else if (X == 9 && Y == 15) begin oled_data = 16'h538c; end
    else if (X == 10 && Y == 15) begin oled_data = 16'h6b4a; end
    else if (X == 13 && Y == 15) begin oled_data = 16'had0f; end
    else if (X == 15 && Y == 15) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 15) begin oled_data = 16'h73af; end
    else if (X == 17 && Y == 15) begin oled_data = 16'had31; end
    else if (X == 18 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 19 && Y == 15) begin oled_data = 16'had31; end
    else if (X == 20 && Y == 15) begin oled_data = 16'had31; end
    else if (X == 21 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 22 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 23 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 24 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 25 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 26 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 27 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 28 && Y == 15) begin oled_data = 16'had31; end
    else if (X == 29 && Y == 15) begin oled_data = 16'had31; end
    else if (X == 30 && Y == 15) begin oled_data = 16'had31; end
    else if (X == 31 && Y == 15) begin oled_data = 16'had31; end
    else if (X >= 32 && X <= 46 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 47 && Y == 15) begin oled_data = 16'h840f; end
    else if (X == 48 && Y == 15) begin oled_data = 16'h840f; end
    else if (X == 49 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 50 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 51 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 52 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 53 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 54 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 55 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 56 && Y == 15) begin oled_data = 16'had31; end
    else if (X == 57 && Y == 15) begin oled_data = 16'had31; end
    else if (X == 58 && Y == 15) begin oled_data = 16'had31; end
    else if (X == 59 && Y == 15) begin oled_data = 16'had31; end
    else if (X == 60 && Y == 15) begin oled_data = 16'had31; end
    else if (X >= 61 && X <= 78 && Y == 15) begin oled_data = 16'ha4f0; end
    else if (X == 79 && Y == 15) begin oled_data = 16'h73af; end
    else if (X == 80 && Y == 15) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 15) begin oled_data = 16'had0f; end
    else if (X == 85 && Y == 15) begin oled_data = 16'hcdd1; end
    else if (X >= 88 && X <= 89 && Y == 15) begin oled_data = 16'h5c27; end
    else if (X == 90 && Y == 15) begin oled_data = 16'h6468; end
    else if (X == 91 && Y == 15) begin oled_data = 16'h64a9; end
    else if (X == 92 && Y == 15) begin oled_data = 16'h64a9; end
    else if (X == 93 && Y == 15) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 15) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 15) begin oled_data = 16'h9551; end
    else if (X == 0 && Y == 16) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 16) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 16) begin oled_data = 16'h4285; end
    else if (X == 3 && Y == 16) begin oled_data = 16'h5b0c; end
    else if (X == 4 && Y == 16) begin oled_data = 16'h8c71; end
    else if (X == 5 && Y == 16) begin oled_data = 16'h538c; end
    else if (X == 6 && Y == 16) begin oled_data = 16'h4b0a; end
    else if (X == 7 && Y == 16) begin oled_data = 16'h5bcd; end
    else if (X == 8 && Y == 16) begin oled_data = 16'h5bcd; end
    else if (X == 9 && Y == 16) begin oled_data = 16'h5bcd; end
    else if (X == 10 && Y == 16) begin oled_data = 16'h83cc; end
    else if (X == 13 && Y == 16) begin oled_data = 16'hb550; end
    else if (X == 15 && Y == 16) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 16) begin oled_data = 16'h840f; end
    else if (X >= 36 && X <= 42 && Y == 16) begin oled_data = 16'hcdd1; end
    else if (X == 47 && Y == 16) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 16) begin oled_data = 16'had31; end
    else if (X >= 71 && X <= 72 && Y == 16) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 16) begin oled_data = 16'h840f; end
    else if (X == 82 && Y == 16) begin oled_data = 16'hb550; end
    else if (X == 88 && Y == 16) begin oled_data = 16'h63e9; end
    else if (X == 89 && Y == 16) begin oled_data = 16'h6468; end
    else if (X == 90 && Y == 16) begin oled_data = 16'h5c27; end
    else if (X == 91 && Y == 16) begin oled_data = 16'h6468; end
    else if (X == 92 && Y == 16) begin oled_data = 16'h64a9; end
    else if (X == 93 && Y == 16) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 16) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 16) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 17) begin oled_data = 16'h9551; end
    else if (X == 1 && Y == 17) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 17) begin oled_data = 16'h4225; end
    else if (X == 3 && Y == 17) begin oled_data = 16'h4a89; end
    else if (X == 4 && Y == 17) begin oled_data = 16'h538c; end
    else if (X == 5 && Y == 17) begin oled_data = 16'h4b0a; end
    else if (X == 6 && Y == 17) begin oled_data = 16'h4b0a; end
    else if (X == 7 && Y == 17) begin oled_data = 16'h5bcd; end
    else if (X == 8 && Y == 17) begin oled_data = 16'h538c; end
    else if (X == 9 && Y == 17) begin oled_data = 16'h6b4a; end
    else if (X == 10 && Y == 17) begin oled_data = 16'h62e8; end
    else if (X == 13 && Y == 17) begin oled_data = 16'hb550; end
    else if (X == 15 && Y == 17) begin oled_data = 16'hbd91; end
    else if (X == 16 && Y == 17) begin oled_data = 16'h840f; end
    else if (X == 18 && Y == 17) begin oled_data = 16'hcdd1; end
    else if (X == 34 && Y == 17) begin oled_data = 16'hbd91; end
    else if (X >= 35 && X <= 36 && Y == 17) begin oled_data = 16'hcdd1; end
    else if (X == 37 && Y == 17) begin oled_data = 16'hbd91; end
    else if (X >= 38 && X <= 44 && Y == 17) begin oled_data = 16'hcdd1; end
    else if (X == 47 && Y == 17) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 17) begin oled_data = 16'had31; end
    else if (X == 56 && Y == 17) begin oled_data = 16'hc5d3; end
    else if (X >= 61 && X <= 74 && Y == 17) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 17) begin oled_data = 16'h8c71; end
    else if (X == 80 && Y == 17) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 17) begin oled_data = 16'had0f; end
    else if (X == 85 && Y == 17) begin oled_data = 16'hcdd1; end
    else if (X == 87 && Y == 17) begin oled_data = 16'hb550; end
    else if (X == 88 && Y == 17) begin oled_data = 16'h63e9; end
    else if (X == 89 && Y == 17) begin oled_data = 16'h6468; end
    else if (X == 90 && Y == 17) begin oled_data = 16'h5c27; end
    else if (X == 91 && Y == 17) begin oled_data = 16'h6468; end
    else if (X == 92 && Y == 17) begin oled_data = 16'h6468; end
    else if (X == 93 && Y == 17) begin oled_data = 16'h64a9; end
    else if (X == 94 && Y == 17) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 17) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 18) begin oled_data = 16'h9551; end
    else if (X == 1 && Y == 18) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 18) begin oled_data = 16'h4225; end
    else if (X == 3 && Y == 18) begin oled_data = 16'h5b0c; end
    else if (X == 4 && Y == 18) begin oled_data = 16'h94b2; end
    else if (X == 5 && Y == 18) begin oled_data = 16'h538c; end
    else if (X == 6 && Y == 18) begin oled_data = 16'h538c; end
    else if (X == 7 && Y == 18) begin oled_data = 16'h5bcd; end
    else if (X == 8 && Y == 18) begin oled_data = 16'h5bcd; end
    else if (X == 9 && Y == 18) begin oled_data = 16'h6b4a; end
    else if (X == 10 && Y == 18) begin oled_data = 16'h62e8; end
    else if (X == 13 && Y == 18) begin oled_data = 16'hb550; end
    else if (X == 15 && Y == 18) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 18) begin oled_data = 16'h840f; end
    else if (X >= 36 && X <= 37 && Y == 18) begin oled_data = 16'hcdd1; end
    else if (X == 47 && Y == 18) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 18) begin oled_data = 16'had31; end
    else if (X == 79 && Y == 18) begin oled_data = 16'h8c71; end
    else if (X == 80 && Y == 18) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 18) begin oled_data = 16'hb550; end
    else if (X == 87 && Y == 18) begin oled_data = 16'h740a; end
    else if (X == 88 && Y == 18) begin oled_data = 16'h5c27; end
    else if (X == 89 && Y == 18) begin oled_data = 16'h6468; end
    else if (X == 90 && Y == 18) begin oled_data = 16'h6468; end
    else if (X == 91 && Y == 18) begin oled_data = 16'h64a9; end
    else if (X == 92 && Y == 18) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 18) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 18) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 18) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 19) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 19) begin oled_data = 16'h53c7; end
    else if (X == 2 && Y == 19) begin oled_data = 16'h4225; end
    else if (X == 3 && Y == 19) begin oled_data = 16'h4a89; end
    else if (X == 4 && Y == 19) begin oled_data = 16'h538c; end
    else if (X == 5 && Y == 19) begin oled_data = 16'h4b0a; end
    else if (X == 6 && Y == 19) begin oled_data = 16'h4b0a; end
    else if (X == 7 && Y == 19) begin oled_data = 16'h538c; end
    else if (X == 8 && Y == 19) begin oled_data = 16'h538c; end
    else if (X == 9 && Y == 19) begin oled_data = 16'h62e8; end
    else if (X == 10 && Y == 19) begin oled_data = 16'h62e8; end
    else if (X == 13 && Y == 19) begin oled_data = 16'had0f; end
    else if (X == 14 && Y == 19) begin oled_data = 16'hcdd1; end
    else if (X == 15 && Y == 19) begin oled_data = 16'hb550; end
    else if (X == 16 && Y == 19) begin oled_data = 16'h840f; end
    else if (X >= 17 && X <= 40 && Y == 19) begin oled_data = 16'hcdd1; end
    else if (X == 47 && Y == 19) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 19) begin oled_data = 16'had31; end
    else if (X >= 53 && X <= 58 && Y == 19) begin oled_data = 16'hcdd1; end
    else if (X == 60 && Y == 19) begin oled_data = 16'hde75; end
    else if (X == 64 && Y == 19) begin oled_data = 16'hcdd1; end
    else if (X == 69 && Y == 19) begin oled_data = 16'hbd91; end
    else if (X >= 70 && X <= 71 && Y == 19) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 19) begin oled_data = 16'h8c71; end
    else if (X >= 80 && X <= 81 && Y == 19) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 19) begin oled_data = 16'had0f; end
    else if (X == 84 && Y == 19) begin oled_data = 16'hb550; end
    else if (X == 85 && Y == 19) begin oled_data = 16'h5b88; end
    else if (X == 86 && Y == 19) begin oled_data = 16'h53c7; end
    else if (X >= 87 && X <= 88 && Y == 19) begin oled_data = 16'h5c27; end
    else if (X == 89 && Y == 19) begin oled_data = 16'h64a9; end
    else if (X == 90 && Y == 19) begin oled_data = 16'h64a9; end
    else if (X == 91 && Y == 19) begin oled_data = 16'h7509; end
    else if (X == 92 && Y == 19) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 19) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 19) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 19) begin oled_data = 16'h9551; end
    else if (X == 0 && Y == 20) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 20) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 20) begin oled_data = 16'h4285; end
    else if (X == 3 && Y == 20) begin oled_data = 16'h5b0c; end
    else if (X == 4 && Y == 20) begin oled_data = 16'h8c71; end
    else if (X == 5 && Y == 20) begin oled_data = 16'h4b0a; end
    else if (X == 6 && Y == 20) begin oled_data = 16'h4b0a; end
    else if (X == 7 && Y == 20) begin oled_data = 16'h5bcd; end
    else if (X == 8 && Y == 20) begin oled_data = 16'h538c; end
    else if (X == 9 && Y == 20) begin oled_data = 16'h62e8; end
    else if (X == 10 && Y == 20) begin oled_data = 16'h62e8; end
    else if (X == 13 && Y == 20) begin oled_data = 16'hb550; end
    else if (X == 15 && Y == 20) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 20) begin oled_data = 16'h840f; end
    else if (X >= 27 && X <= 37 && Y == 20) begin oled_data = 16'hcdd1; end
    else if (X == 47 && Y == 20) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 20) begin oled_data = 16'hb573; end
    else if (X == 56 && Y == 20) begin oled_data = 16'hde75; end
    else if (X == 62 && Y == 20) begin oled_data = 16'hde75; end
    else if (X >= 67 && X <= 69 && Y == 20) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 20) begin oled_data = 16'h8c71; end
    else if (X == 80 && Y == 20) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 20) begin oled_data = 16'hb550; end
    else if (X == 84 && Y == 20) begin oled_data = 16'hb550; end
    else if (X == 85 && Y == 20) begin oled_data = 16'h53c7; end
    else if (X == 86 && Y == 20) begin oled_data = 16'h5c27; end
    else if (X == 87 && Y == 20) begin oled_data = 16'h6468; end
    else if (X == 88 && Y == 20) begin oled_data = 16'h6468; end
    else if (X == 89 && Y == 20) begin oled_data = 16'h7509; end
    else if (X == 90 && Y == 20) begin oled_data = 16'h7509; end
    else if (X == 91 && Y == 20) begin oled_data = 16'h7d6b; end
    else if (X == 92 && Y == 20) begin oled_data = 16'h7d6b; end
    else if (X == 93 && Y == 20) begin oled_data = 16'h7d6b; end
    else if (X == 94 && Y == 20) begin oled_data = 16'h7509; end
    else if (X == 95 && Y == 20) begin oled_data = 16'h8d0f; end
    else if (X == 0 && Y == 21) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 21) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 21) begin oled_data = 16'h4285; end
    else if (X == 3 && Y == 21) begin oled_data = 16'h4a27; end
    else if (X == 4 && Y == 21) begin oled_data = 16'h4a89; end
    else if (X == 5 && Y == 21) begin oled_data = 16'h4a27; end
    else if (X == 6 && Y == 21) begin oled_data = 16'h4a27; end
    else if (X == 7 && Y == 21) begin oled_data = 16'h4a89; end
    else if (X == 8 && Y == 21) begin oled_data = 16'h4a89; end
    else if (X == 9 && Y == 21) begin oled_data = 16'h5a87; end
    else if (X == 10 && Y == 21) begin oled_data = 16'h5a87; end
    else if (X == 13 && Y == 21) begin oled_data = 16'hb550; end
    else if (X == 15 && Y == 21) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 21) begin oled_data = 16'h840f; end
    else if (X == 21 && Y == 21) begin oled_data = 16'hde75; end
    else if (X == 23 && Y == 21) begin oled_data = 16'hde75; end
    else if (X == 30 && Y == 21) begin oled_data = 16'hcdd1; end
    else if (X == 33 && Y == 21) begin oled_data = 16'hde75; end
    else if (X == 37 && Y == 21) begin oled_data = 16'hcdd1; end
    else if (X == 44 && Y == 21) begin oled_data = 16'hde75; end
    else if (X == 47 && Y == 21) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 21) begin oled_data = 16'had31; end
    else if (X == 54 && Y == 21) begin oled_data = 16'hde75; end
    else if (X == 61 && Y == 21) begin oled_data = 16'hde75; end
    else if (X == 64 && Y == 21) begin oled_data = 16'hde75; end
    else if (X == 71 && Y == 21) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 21) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 21) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 21) begin oled_data = 16'had0f; end
    else if (X == 84 && Y == 21) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 21) begin oled_data = 16'h53c7; end
    else if (X == 86 && Y == 21) begin oled_data = 16'h5c27; end
    else if (X == 87 && Y == 21) begin oled_data = 16'h6468; end
    else if (X == 88 && Y == 21) begin oled_data = 16'h64a9; end
    else if (X == 89 && Y == 21) begin oled_data = 16'h7509; end
    else if (X == 90 && Y == 21) begin oled_data = 16'h7d6b; end
    else if (X == 91 && Y == 21) begin oled_data = 16'h7d6b; end
    else if (X == 92 && Y == 21) begin oled_data = 16'h7d6b; end
    else if (X == 93 && Y == 21) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 21) begin oled_data = 16'h7509; end
    else if (X == 95 && Y == 21) begin oled_data = 16'h8d0f; end
    else if (X == 0 && Y == 22) begin oled_data = 16'hb5b6; end
    else if (X == 1 && Y == 22) begin oled_data = 16'h848c; end
    else if (X == 2 && Y == 22) begin oled_data = 16'h83cc; end
    else if (X == 3 && Y == 22) begin oled_data = 16'h83cc; end
    else if (X == 4 && Y == 22) begin oled_data = 16'h83cc; end
    else if (X == 5 && Y == 22) begin oled_data = 16'h940c; end
    else if (X == 6 && Y == 22) begin oled_data = 16'h940c; end
    else if (X == 7 && Y == 22) begin oled_data = 16'h940c; end
    else if (X == 8 && Y == 22) begin oled_data = 16'h940c; end
    else if (X == 9 && Y == 22) begin oled_data = 16'h940c; end
    else if (X == 10 && Y == 22) begin oled_data = 16'h940c; end
    else if (X == 13 && Y == 22) begin oled_data = 16'had0f; end
    else if (X == 15 && Y == 22) begin oled_data = 16'hbd91; end
    else if (X == 16 && Y == 22) begin oled_data = 16'h840f; end
    else if (X >= 17 && X <= 34 && Y == 22) begin oled_data = 16'hcdd1; end
    else if (X == 45 && Y == 22) begin oled_data = 16'hc5d3; end
    else if (X == 47 && Y == 22) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 22) begin oled_data = 16'had31; end
    else if (X == 55 && Y == 22) begin oled_data = 16'hcdd1; end
    else if (X == 58 && Y == 22) begin oled_data = 16'hde75; end
    else if (X == 69 && Y == 22) begin oled_data = 16'hbd91; end
    else if (X >= 71 && X <= 77 && Y == 22) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 22) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 22) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 22) begin oled_data = 16'ha4f0; end
    else if (X >= 83 && X <= 84 && Y == 22) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 22) begin oled_data = 16'h63e9; end
    else if (X == 86 && Y == 22) begin oled_data = 16'h5c27; end
    else if (X == 87 && Y == 22) begin oled_data = 16'h6468; end
    else if (X == 88 && Y == 22) begin oled_data = 16'h64a9; end
    else if (X == 89 && Y == 22) begin oled_data = 16'h7509; end
    else if (X == 90 && Y == 22) begin oled_data = 16'h7509; end
    else if (X == 91 && Y == 22) begin oled_data = 16'h7509; end
    else if (X == 92 && Y == 22) begin oled_data = 16'h7d6b; end
    else if (X == 93 && Y == 22) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 22) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 22) begin oled_data = 16'h8d0f; end
    else if (X == 0 && Y == 23) begin oled_data = 16'hce16; end
    else if (X == 5 && Y == 23) begin oled_data = 16'hcdd1; end
    else if (X == 13 && Y == 23) begin oled_data = 16'hb550; end
    else if (X == 15 && Y == 23) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 23) begin oled_data = 16'h840f; end
    else if (X >= 32 && X <= 36 && Y == 23) begin oled_data = 16'hcdd1; end
    else if (X == 47 && Y == 23) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 23) begin oled_data = 16'had31; end
    else if (X == 51 && Y == 23) begin oled_data = 16'hde75; end
    else if (X == 67 && Y == 23) begin oled_data = 16'hde75; end
    else if (X == 79 && Y == 23) begin oled_data = 16'h8c71; end
    else if (X == 82 && Y == 23) begin oled_data = 16'hb550; end
    else if (X == 85 && Y == 23) begin oled_data = 16'h740a; end
    else if (X == 86 && Y == 23) begin oled_data = 16'h5c27; end
    else if (X == 87 && Y == 23) begin oled_data = 16'h64a9; end
    else if (X == 88 && Y == 23) begin oled_data = 16'h64a9; end
    else if (X == 89 && Y == 23) begin oled_data = 16'h7509; end
    else if (X == 90 && Y == 23) begin oled_data = 16'h7509; end
    else if (X == 91 && Y == 23) begin oled_data = 16'h7d6b; end
    else if (X == 92 && Y == 23) begin oled_data = 16'h7d6b; end
    else if (X == 93 && Y == 23) begin oled_data = 16'h7d6b; end
    else if (X == 94 && Y == 23) begin oled_data = 16'h7d6b; end
    else if (X == 95 && Y == 23) begin oled_data = 16'h8d0f; end
    else if (X == 0 && Y == 24) begin oled_data = 16'hce16; end
    else if (X == 2 && Y == 24) begin oled_data = 16'hcdd1; end
    else if (X == 4 && Y == 24) begin oled_data = 16'had0f; end
    else if (X == 5 && Y == 24) begin oled_data = 16'h4b07; end
    else if (X == 7 && Y == 24) begin oled_data = 16'hb550; end
    else if (X == 8 && Y == 24) begin oled_data = 16'had0f; end
    else if (X == 9 && Y == 24) begin oled_data = 16'hbd91; end
    else if (X == 10 && Y == 24) begin oled_data = 16'had0f; end
    else if (X == 11 && Y == 24) begin oled_data = 16'hbd91; end
    else if (X == 12 && Y == 24) begin oled_data = 16'hbd91; end
    else if (X == 13 && Y == 24) begin oled_data = 16'h9c8e; end
    else if (X == 15 && Y == 24) begin oled_data = 16'hb550; end
    else if (X == 16 && Y == 24) begin oled_data = 16'h840f; end
    else if (X == 20 && Y == 24) begin oled_data = 16'hde75; end
    else if (X >= 24 && X <= 28 && Y == 24) begin oled_data = 16'hcdd1; end
    else if (X == 29 && Y == 24) begin oled_data = 16'hbd91; end
    else if (X >= 32 && X <= 38 && Y == 24) begin oled_data = 16'hcdd1; end
    else if (X == 44 && Y == 24) begin oled_data = 16'hbd91; end
    else if (X == 45 && Y == 24) begin oled_data = 16'had31; end
    else if (X == 46 && Y == 24) begin oled_data = 16'had31; end
    else if (X == 47 && Y == 24) begin oled_data = 16'h8c71; end
    else if (X == 48 && Y == 24) begin oled_data = 16'h8c71; end
    else if (X == 49 && Y == 24) begin oled_data = 16'had31; end
    else if (X == 50 && Y == 24) begin oled_data = 16'had31; end
    else if (X >= 51 && X <= 75 && Y == 24) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 24) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 24) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 24) begin oled_data = 16'h9c8e; end
    else if (X == 84 && Y == 24) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 24) begin oled_data = 16'h63e9; end
    else if (X == 86 && Y == 24) begin oled_data = 16'h6468; end
    else if (X == 87 && Y == 24) begin oled_data = 16'h6468; end
    else if (X == 88 && Y == 24) begin oled_data = 16'h6468; end
    else if (X == 89 && Y == 24) begin oled_data = 16'h6468; end
    else if (X == 90 && Y == 24) begin oled_data = 16'h7509; end
    else if (X == 91 && Y == 24) begin oled_data = 16'h7d6b; end
    else if (X == 92 && Y == 24) begin oled_data = 16'h7d6b; end
    else if (X == 93 && Y == 24) begin oled_data = 16'h7d6b; end
    else if (X == 94 && Y == 24) begin oled_data = 16'h7509; end
    else if (X == 95 && Y == 24) begin oled_data = 16'h8d0f; end
    else if (X == 0 && Y == 25) begin oled_data = 16'hce16; end
    else if (X == 4 && Y == 25) begin oled_data = 16'hb550; end
    else if (X == 5 && Y == 25) begin oled_data = 16'h5b88; end
    else if (X >= 6 && X <= 15 && Y == 25) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 25) begin oled_data = 16'h840f; end
    else if (X >= 26 && X <= 39 && Y == 25) begin oled_data = 16'hcdd1; end
    else if (X == 42 && Y == 25) begin oled_data = 16'had31; end
    else if (X == 43 && Y == 25) begin oled_data = 16'h8c71; end
    else if (X == 44 && Y == 25) begin oled_data = 16'h8c71; end
    else if (X == 45 && Y == 25) begin oled_data = 16'ha4f0; end
    else if (X == 46 && Y == 25) begin oled_data = 16'hbd72; end
    else if (X == 47 && Y == 25) begin oled_data = 16'ha4f0; end
    else if (X == 48 && Y == 25) begin oled_data = 16'h9cb1; end
    else if (X == 49 && Y == 25) begin oled_data = 16'had31; end
    else if (X == 50 && Y == 25) begin oled_data = 16'h9cb1; end
    else if (X == 51 && Y == 25) begin oled_data = 16'h8c71; end
    else if (X == 52 && Y == 25) begin oled_data = 16'h840f; end
    else if (X == 53 && Y == 25) begin oled_data = 16'had31; end
    else if (X == 73 && Y == 25) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 25) begin oled_data = 16'h840f; end
    else if (X >= 80 && X <= 84 && Y == 25) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 25) begin oled_data = 16'h53c7; end
    else if (X >= 86 && X <= 87 && Y == 25) begin oled_data = 16'h5c27; end
    else if (X == 88 && Y == 25) begin oled_data = 16'h6468; end
    else if (X == 89 && Y == 25) begin oled_data = 16'h64a9; end
    else if (X == 90 && Y == 25) begin oled_data = 16'h64a9; end
    else if (X == 91 && Y == 25) begin oled_data = 16'h7509; end
    else if (X == 92 && Y == 25) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 25) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 25) begin oled_data = 16'h7509; end
    else if (X == 95 && Y == 25) begin oled_data = 16'h8d0f; end
    else if (X == 0 && Y == 26) begin oled_data = 16'hce16; end
    else if (X == 3 && Y == 26) begin oled_data = 16'hcdd1; end
    else if (X == 4 && Y == 26) begin oled_data = 16'h740a; end
    else if (X == 5 && Y == 26) begin oled_data = 16'h4b07; end
    else if (X == 6 && Y == 26) begin oled_data = 16'h948d; end
    else if (X == 7 && Y == 26) begin oled_data = 16'ha4ee; end
    else if (X == 8 && Y == 26) begin oled_data = 16'ha4ee; end
    else if (X == 9 && Y == 26) begin oled_data = 16'had0f; end
    else if (X == 10 && Y == 26) begin oled_data = 16'h9cad; end
    else if (X == 11 && Y == 26) begin oled_data = 16'h948d; end
    else if (X == 12 && Y == 26) begin oled_data = 16'ha4ee; end
    else if (X == 13 && Y == 26) begin oled_data = 16'h948d; end
    else if (X >= 14 && X <= 15 && Y == 26) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 26) begin oled_data = 16'h840f; end
    else if (X == 20 && Y == 26) begin oled_data = 16'hde75; end
    else if (X == 23 && Y == 26) begin oled_data = 16'hde75; end
    else if (X == 32 && Y == 26) begin oled_data = 16'hde75; end
    else if (X == 35 && Y == 26) begin oled_data = 16'hde75; end
    else if (X == 40 && Y == 26) begin oled_data = 16'had31; end
    else if (X == 41 && Y == 26) begin oled_data = 16'h8c71; end
    else if (X == 42 && Y == 26) begin oled_data = 16'had31; end
    else if (X == 47 && Y == 26) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 26) begin oled_data = 16'had31; end
    else if (X >= 50 && X <= 52 && Y == 26) begin oled_data = 16'hcdd1; end
    else if (X == 53 && Y == 26) begin oled_data = 16'ha4f0; end
    else if (X == 54 && Y == 26) begin oled_data = 16'h840f; end
    else if (X == 55 && Y == 26) begin oled_data = 16'ha4f0; end
    else if (X == 60 && Y == 26) begin oled_data = 16'hde75; end
    else if (X == 63 && Y == 26) begin oled_data = 16'hde75; end
    else if (X == 64 && Y == 26) begin oled_data = 16'hde75; end
    else if (X == 68 && Y == 26) begin oled_data = 16'hde75; end
    else if (X == 72 && Y == 26) begin oled_data = 16'hde75; end
    else if (X == 74 && Y == 26) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 26) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 26) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 26) begin oled_data = 16'hbd91; end
    else if (X == 84 && Y == 26) begin oled_data = 16'hbd91; end
    else if (X == 85 && Y == 26) begin oled_data = 16'h4b07; end
    else if (X == 86 && Y == 26) begin oled_data = 16'h53c7; end
    else if (X == 87 && Y == 26) begin oled_data = 16'h53c7; end
    else if (X == 88 && Y == 26) begin oled_data = 16'h5c27; end
    else if (X == 89 && Y == 26) begin oled_data = 16'h6468; end
    else if (X == 90 && Y == 26) begin oled_data = 16'h5bc8; end
    else if (X == 91 && Y == 26) begin oled_data = 16'h6468; end
    else if (X == 92 && Y == 26) begin oled_data = 16'h64a9; end
    else if (X == 93 && Y == 26) begin oled_data = 16'h64a9; end
    else if (X == 94 && Y == 26) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 26) begin oled_data = 16'h8d0f; end
    else if (X == 0 && Y == 27) begin oled_data = 16'hb573; end
    else if (X == 1 && Y == 27) begin oled_data = 16'h740a; end
    else if (X == 2 && Y == 27) begin oled_data = 16'h53c7; end
    else if (X >= 3 && X <= 4 && Y == 27) begin oled_data = 16'h5c27; end
    else if (X == 5 && Y == 27) begin oled_data = 16'h4b07; end
    else if (X == 6 && Y == 27) begin oled_data = 16'h53c7; end
    else if (X == 7 && Y == 27) begin oled_data = 16'h53c7; end
    else if (X == 8 && Y == 27) begin oled_data = 16'h4346; end
    else if (X == 9 && Y == 27) begin oled_data = 16'h53c7; end
    else if (X == 10 && Y == 27) begin oled_data = 16'h4346; end
    else if (X == 11 && Y == 27) begin oled_data = 16'h53c7; end
    else if (X == 12 && Y == 27) begin oled_data = 16'h53c7; end
    else if (X == 13 && Y == 27) begin oled_data = 16'h53c7; end
    else if (X == 14 && Y == 27) begin oled_data = 16'h740a; end
    else if (X == 15 && Y == 27) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 27) begin oled_data = 16'h840f; end
    else if (X >= 17 && X <= 30 && Y == 27) begin oled_data = 16'hcdd1; end
    else if (X == 34 && Y == 27) begin oled_data = 16'hc5b2; end
    else if (X == 37 && Y == 27) begin oled_data = 16'hde75; end
    else if (X == 39 && Y == 27) begin oled_data = 16'h94b2; end
    else if (X == 40 && Y == 27) begin oled_data = 16'had31; end
    else if (X == 45 && Y == 27) begin oled_data = 16'hbd91; end
    else if (X == 47 && Y == 27) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 27) begin oled_data = 16'ha4f0; end
    else if (X >= 49 && X <= 54 && Y == 27) begin oled_data = 16'hcdd1; end
    else if (X == 55 && Y == 27) begin oled_data = 16'h9cb1; end
    else if (X == 56 && Y == 27) begin oled_data = 16'h840f; end
    else if (X >= 58 && X <= 59 && Y == 27) begin oled_data = 16'hcdd1; end
    else if (X == 66 && Y == 27) begin oled_data = 16'hc5b2; end
    else if (X >= 69 && X <= 74 && Y == 27) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 27) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 27) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 27) begin oled_data = 16'ha4f0; end
    else if (X == 83 && Y == 27) begin oled_data = 16'hbd91; end
    else if (X == 84 && Y == 27) begin oled_data = 16'hbd91; end
    else if (X == 85 && Y == 27) begin oled_data = 16'h948d; end
    else if (X == 86 && Y == 27) begin oled_data = 16'h740a; end
    else if (X == 87 && Y == 27) begin oled_data = 16'h740a; end
    else if (X == 88 && Y == 27) begin oled_data = 16'h5b88; end
    else if (X == 89 && Y == 27) begin oled_data = 16'h4346; end
    else if (X == 90 && Y == 27) begin oled_data = 16'h4b07; end
    else if (X == 91 && Y == 27) begin oled_data = 16'h5c27; end
    else if (X == 92 && Y == 27) begin oled_data = 16'h6468; end
    else if (X == 93 && Y == 27) begin oled_data = 16'h64a9; end
    else if (X == 94 && Y == 27) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 27) begin oled_data = 16'h8d0f; end
    else if (X == 0 && Y == 28) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 28) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 28) begin oled_data = 16'h6468; end
    else if (X == 3 && Y == 28) begin oled_data = 16'h5c27; end
    else if (X == 4 && Y == 28) begin oled_data = 16'h6468; end
    else if (X == 5 && Y == 28) begin oled_data = 16'h53c7; end
    else if (X == 6 && Y == 28) begin oled_data = 16'h5c27; end
    else if (X == 7 && Y == 28) begin oled_data = 16'h53c7; end
    else if (X == 8 && Y == 28) begin oled_data = 16'h53c7; end
    else if (X == 9 && Y == 28) begin oled_data = 16'h5c27; end
    else if (X == 10 && Y == 28) begin oled_data = 16'h53c7; end
    else if (X >= 11 && X <= 12 && Y == 28) begin oled_data = 16'h5c27; end
    else if (X == 13 && Y == 28) begin oled_data = 16'h740a; end
    else if (X == 14 && Y == 28) begin oled_data = 16'had0f; end
    else if (X == 15 && Y == 28) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 28) begin oled_data = 16'h840f; end
    else if (X >= 21 && X <= 24 && Y == 28) begin oled_data = 16'hcdd1; end
    else if (X == 36 && Y == 28) begin oled_data = 16'hde75; end
    else if (X == 37 && Y == 28) begin oled_data = 16'hc5d3; end
    else if (X == 38 && Y == 28) begin oled_data = 16'h94b2; end
    else if (X == 39 && Y == 28) begin oled_data = 16'hc5d4; end
    else if (X == 41 && Y == 28) begin oled_data = 16'hde75; end
    else if (X == 42 && Y == 28) begin oled_data = 16'hde75; end
    else if (X == 45 && Y == 28) begin oled_data = 16'hde75; end
    else if (X == 47 && Y == 28) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 28) begin oled_data = 16'had31; end
    else if (X >= 50 && X <= 53 && Y == 28) begin oled_data = 16'hcdd1; end
    else if (X == 56 && Y == 28) begin oled_data = 16'hb550; end
    else if (X == 57 && Y == 28) begin oled_data = 16'h840f; end
    else if (X == 79 && Y == 28) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 28) begin oled_data = 16'hcdd1; end
    else if (X == 89 && Y == 28) begin oled_data = 16'h848c; end
    else if (X == 90 && Y == 28) begin oled_data = 16'h4346; end
    else if (X == 91 && Y == 28) begin oled_data = 16'h5c27; end
    else if (X == 92 && Y == 28) begin oled_data = 16'h6468; end
    else if (X == 93 && Y == 28) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 28) begin oled_data = 16'h7509; end
    else if (X == 95 && Y == 28) begin oled_data = 16'h8d0f; end
    else if (X == 0 && Y == 29) begin oled_data = 16'ha593; end
    else if (X >= 1 && X <= 2 && Y == 29) begin oled_data = 16'h5c27; end
    else if (X == 3 && Y == 29) begin oled_data = 16'h6468; end
    else if (X == 4 && Y == 29) begin oled_data = 16'h5c27; end
    else if (X == 5 && Y == 29) begin oled_data = 16'h4346; end
    else if (X == 6 && Y == 29) begin oled_data = 16'h53c7; end
    else if (X == 7 && Y == 29) begin oled_data = 16'h53c7; end
    else if (X == 8 && Y == 29) begin oled_data = 16'h63e9; end
    else if (X == 9 && Y == 29) begin oled_data = 16'h53c7; end
    else if (X == 10 && Y == 29) begin oled_data = 16'h53c7; end
    else if (X == 11 && Y == 29) begin oled_data = 16'h848c; end
    else if (X == 12 && Y == 29) begin oled_data = 16'hb550; end
    else if (X == 13 && Y == 29) begin oled_data = 16'had0f; end
    else if (X == 14 && Y == 29) begin oled_data = 16'h9cb1; end
    else if (X == 15 && Y == 29) begin oled_data = 16'h840f; end
    else if (X == 16 && Y == 29) begin oled_data = 16'h840f; end
    else if (X >= 17 && X <= 20 && Y == 29) begin oled_data = 16'hcdd1; end
    else if (X == 21 && Y == 29) begin oled_data = 16'hbd91; end
    else if (X >= 22 && X <= 26 && Y == 29) begin oled_data = 16'hcdd1; end
    else if (X == 30 && Y == 29) begin oled_data = 16'hde75; end
    else if (X == 33 && Y == 29) begin oled_data = 16'hde75; end
    else if (X == 37 && Y == 29) begin oled_data = 16'h94b2; end
    else if (X == 38 && Y == 29) begin oled_data = 16'hc5d4; end
    else if (X == 39 && Y == 29) begin oled_data = 16'hde75; end
    else if (X == 40 && Y == 29) begin oled_data = 16'hde75; end
    else if (X == 41 && Y == 29) begin oled_data = 16'hde75; end
    else if (X == 45 && Y == 29) begin oled_data = 16'hc5b2; end
    else if (X == 47 && Y == 29) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 29) begin oled_data = 16'ha4f0; end
    else if (X >= 49 && X <= 50 && Y == 29) begin oled_data = 16'hcdd1; end
    else if (X == 53 && Y == 29) begin oled_data = 16'hb550; end
    else if (X >= 54 && X <= 56 && Y == 29) begin oled_data = 16'hcdd1; end
    else if (X == 57 && Y == 29) begin oled_data = 16'hb550; end
    else if (X == 58 && Y == 29) begin oled_data = 16'h840f; end
    else if (X == 60 && Y == 29) begin oled_data = 16'hde75; end
    else if (X == 70 && Y == 29) begin oled_data = 16'hcdd1; end
    else if (X == 74 && Y == 29) begin oled_data = 16'hbd91; end
    else if (X == 77 && Y == 29) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 29) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 29) begin oled_data = 16'h840f; end
    else if (X == 81 && Y == 29) begin oled_data = 16'h9cb1; end
    else if (X == 82 && Y == 29) begin oled_data = 16'ha4f0; end
    else if (X == 90 && Y == 29) begin oled_data = 16'h5b88; end
    else if (X == 91 && Y == 29) begin oled_data = 16'h5c27; end
    else if (X == 92 && Y == 29) begin oled_data = 16'h64a9; end
    else if (X == 93 && Y == 29) begin oled_data = 16'h64a9; end
    else if (X == 94 && Y == 29) begin oled_data = 16'h7509; end
    else if (X == 95 && Y == 29) begin oled_data = 16'h8d0f; end
    else if (X == 0 && Y == 30) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 30) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 30) begin oled_data = 16'h53c7; end
    else if (X == 3 && Y == 30) begin oled_data = 16'h6468; end
    else if (X == 4 && Y == 30) begin oled_data = 16'h6468; end
    else if (X == 5 && Y == 30) begin oled_data = 16'h53c7; end
    else if (X == 6 && Y == 30) begin oled_data = 16'h9cad; end
    else if (X == 7 && Y == 30) begin oled_data = 16'h7c4b; end
    else if (X == 8 && Y == 30) begin oled_data = 16'h53c7; end
    else if (X == 9 && Y == 30) begin oled_data = 16'h740a; end
    else if (X == 10 && Y == 30) begin oled_data = 16'hbd91; end
    else if (X == 11 && Y == 30) begin oled_data = 16'had31; end
    else if (X == 12 && Y == 30) begin oled_data = 16'h840f; end
    else if (X == 13 && Y == 30) begin oled_data = 16'h840d; end
    else if (X == 14 && Y == 30) begin oled_data = 16'had0f; end
    else if (X == 15 && Y == 30) begin oled_data = 16'hb550; end
    else if (X == 16 && Y == 30) begin oled_data = 16'h840d; end
    else if (X >= 17 && X <= 23 && Y == 30) begin oled_data = 16'hcdd1; end
    else if (X == 36 && Y == 30) begin oled_data = 16'ha514; end
    else if (X == 37 && Y == 30) begin oled_data = 16'had31; end
    else if (X == 38 && Y == 30) begin oled_data = 16'hde75; end
    else if (X == 39 && Y == 30) begin oled_data = 16'hde75; end
    else if (X == 40 && Y == 30) begin oled_data = 16'hde75; end
    else if (X == 41 && Y == 30) begin oled_data = 16'hde75; end
    else if (X == 42 && Y == 30) begin oled_data = 16'hde75; end
    else if (X == 43 && Y == 30) begin oled_data = 16'hde75; end
    else if (X == 44 && Y == 30) begin oled_data = 16'hde75; end
    else if (X == 45 && Y == 30) begin oled_data = 16'hde75; end
    else if (X == 46 && Y == 30) begin oled_data = 16'hde75; end
    else if (X == 47 && Y == 30) begin oled_data = 16'hb573; end
    else if (X == 48 && Y == 30) begin oled_data = 16'had31; end
    else if (X >= 50 && X <= 53 && Y == 30) begin oled_data = 16'hcdd1; end
    else if (X == 58 && Y == 30) begin oled_data = 16'ha4f0; end
    else if (X == 59 && Y == 30) begin oled_data = 16'h9cb1; end
    else if (X == 78 && Y == 30) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 30) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 30) begin oled_data = 16'hb550; end
    else if (X == 81 && Y == 30) begin oled_data = 16'had31; end
    else if (X == 82 && Y == 30) begin oled_data = 16'h8c71; end
    else if (X == 83 && Y == 30) begin oled_data = 16'h8c71; end
    else if (X == 84 && Y == 30) begin oled_data = 16'hbd72; end
    else if (X == 86 && Y == 30) begin oled_data = 16'hde75; end
    else if (X == 90 && Y == 30) begin oled_data = 16'h948d; end
    else if (X == 91 && Y == 30) begin oled_data = 16'h5c27; end
    else if (X == 92 && Y == 30) begin oled_data = 16'h64a9; end
    else if (X == 93 && Y == 30) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 30) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 30) begin oled_data = 16'h84ce; end
    else if (X == 0 && Y == 31) begin oled_data = 16'ha593; end
    else if (X >= 1 && X <= 2 && Y == 31) begin oled_data = 16'h5c27; end
    else if (X == 3 && Y == 31) begin oled_data = 16'h6468; end
    else if (X == 4 && Y == 31) begin oled_data = 16'h64a9; end
    else if (X == 5 && Y == 31) begin oled_data = 16'h5c27; end
    else if (X == 6 && Y == 31) begin oled_data = 16'h948d; end
    else if (X == 7 && Y == 31) begin oled_data = 16'h5bc8; end
    else if (X == 8 && Y == 31) begin oled_data = 16'h5bc8; end
    else if (X == 9 && Y == 31) begin oled_data = 16'hb550; end
    else if (X == 10 && Y == 31) begin oled_data = 16'h8c71; end
    else if (X == 11 && Y == 31) begin oled_data = 16'h8c71; end
    else if (X >= 12 && X <= 15 && Y == 31) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 31) begin oled_data = 16'h840f; end
    else if (X >= 17 && X <= 27 && Y == 31) begin oled_data = 16'hcdd1; end
    else if (X == 35 && Y == 31) begin oled_data = 16'hc5d3; end
    else if (X == 36 && Y == 31) begin oled_data = 16'h8c71; end
    else if (X == 39 && Y == 31) begin oled_data = 16'hde75; end
    else if (X == 42 && Y == 31) begin oled_data = 16'hde75; end
    else if (X == 43 && Y == 31) begin oled_data = 16'hde75; end
    else if (X == 44 && Y == 31) begin oled_data = 16'hde75; end
    else if (X == 45 && Y == 31) begin oled_data = 16'hde75; end
    else if (X == 46 && Y == 31) begin oled_data = 16'hde75; end
    else if (X == 47 && Y == 31) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 31) begin oled_data = 16'had31; end
    else if (X >= 49 && X <= 58 && Y == 31) begin oled_data = 16'hcdd1; end
    else if (X == 59 && Y == 31) begin oled_data = 16'h840f; end
    else if (X == 60 && Y == 31) begin oled_data = 16'hcdd1; end
    else if (X == 65 && Y == 31) begin oled_data = 16'hde75; end
    else if (X == 67 && Y == 31) begin oled_data = 16'hde75; end
    else if (X >= 77 && X <= 78 && Y == 31) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 31) begin oled_data = 16'h840f; end
    else if (X >= 80 && X <= 83 && Y == 31) begin oled_data = 16'hcdd1; end
    else if (X == 84 && Y == 31) begin oled_data = 16'h8c71; end
    else if (X == 85 && Y == 31) begin oled_data = 16'h8c71; end
    else if (X == 90 && Y == 31) begin oled_data = 16'ha4f0; end
    else if (X == 91 && Y == 31) begin oled_data = 16'h5c27; end
    else if (X == 92 && Y == 31) begin oled_data = 16'h64a9; end
    else if (X == 93 && Y == 31) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 31) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 31) begin oled_data = 16'h84ce; end
    else if (X == 0 && Y == 32) begin oled_data = 16'h9551; end
    else if (X == 1 && Y == 32) begin oled_data = 16'h6468; end
    else if (X == 2 && Y == 32) begin oled_data = 16'h6468; end
    else if (X == 3 && Y == 32) begin oled_data = 16'h64a9; end
    else if (X == 4 && Y == 32) begin oled_data = 16'h64a9; end
    else if (X >= 5 && X <= 7 && Y == 32) begin oled_data = 16'h5c27; end
    else if (X == 8 && Y == 32) begin oled_data = 16'ha4ee; end
    else if (X == 9 && Y == 32) begin oled_data = 16'h8c71; end
    else if (X == 10 && Y == 32) begin oled_data = 16'ha4f0; end
    else if (X >= 13 && X <= 15 && Y == 32) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 32) begin oled_data = 16'h840f; end
    else if (X >= 17 && X <= 29 && Y == 32) begin oled_data = 16'hcdd1; end
    else if (X == 35 && Y == 32) begin oled_data = 16'h94b2; end
    else if (X == 36 && Y == 32) begin oled_data = 16'hc5d3; end
    else if (X == 43 && Y == 32) begin oled_data = 16'hde75; end
    else if (X == 44 && Y == 32) begin oled_data = 16'hde75; end
    else if (X == 45 && Y == 32) begin oled_data = 16'hde75; end
    else if (X == 47 && Y == 32) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 32) begin oled_data = 16'ha4f0; end
    else if (X >= 49 && X <= 58 && Y == 32) begin oled_data = 16'hcdd1; end
    else if (X == 59 && Y == 32) begin oled_data = 16'hb550; end
    else if (X == 60 && Y == 32) begin oled_data = 16'h9cb1; end
    else if (X >= 75 && X <= 77 && Y == 32) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 32) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 32) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 32) begin oled_data = 16'h9cb1; end
    else if (X == 86 && Y == 32) begin oled_data = 16'h9cb1; end
    else if (X == 90 && Y == 32) begin oled_data = 16'h740a; end
    else if (X == 91 && Y == 32) begin oled_data = 16'h5c27; end
    else if (X == 92 && Y == 32) begin oled_data = 16'h6468; end
    else if (X == 93 && Y == 32) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 32) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 32) begin oled_data = 16'h8d0f; end
    else if (X == 0 && Y == 33) begin oled_data = 16'h9551; end
    else if (X == 1 && Y == 33) begin oled_data = 16'h64a9; end
    else if (X == 2 && Y == 33) begin oled_data = 16'h64a9; end
    else if (X == 3 && Y == 33) begin oled_data = 16'h64a9; end
    else if (X == 4 && Y == 33) begin oled_data = 16'h64a9; end
    else if (X >= 5 && X <= 6 && Y == 33) begin oled_data = 16'h5c27; end
    else if (X == 7 && Y == 33) begin oled_data = 16'h740a; end
    else if (X == 8 && Y == 33) begin oled_data = 16'hbd91; end
    else if (X == 9 && Y == 33) begin oled_data = 16'h8c71; end
    else if (X >= 10 && X <= 15 && Y == 33) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 33) begin oled_data = 16'h840f; end
    else if (X == 27 && Y == 33) begin oled_data = 16'hcdd1; end
    else if (X == 35 && Y == 33) begin oled_data = 16'h8c71; end
    else if (X == 47 && Y == 33) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 33) begin oled_data = 16'had31; end
    else if (X >= 50 && X <= 58 && Y == 33) begin oled_data = 16'hcdd1; end
    else if (X == 60 && Y == 33) begin oled_data = 16'h840f; end
    else if (X >= 74 && X <= 77 && Y == 33) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 33) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 33) begin oled_data = 16'hcdd1; end
    else if (X == 86 && Y == 33) begin oled_data = 16'h840f; end
    else if (X == 87 && Y == 33) begin oled_data = 16'hbd91; end
    else if (X == 90 && Y == 33) begin oled_data = 16'h63e9; end
    else if (X >= 91 && X <= 92 && Y == 33) begin oled_data = 16'h5c27; end
    else if (X == 93 && Y == 33) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 33) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 33) begin oled_data = 16'h9551; end
    else if (X == 0 && Y == 34) begin oled_data = 16'h9551; end
    else if (X == 1 && Y == 34) begin oled_data = 16'h64a9; end
    else if (X == 2 && Y == 34) begin oled_data = 16'h5c27; end
    else if (X == 3 && Y == 34) begin oled_data = 16'h6468; end
    else if (X == 4 && Y == 34) begin oled_data = 16'h64a9; end
    else if (X == 5 && Y == 34) begin oled_data = 16'h53c7; end
    else if (X == 6 && Y == 34) begin oled_data = 16'h53c7; end
    else if (X == 7 && Y == 34) begin oled_data = 16'had0f; end
    else if (X == 8 && Y == 34) begin oled_data = 16'h840f; end
    else if (X == 9 && Y == 34) begin oled_data = 16'hbd91; end
    else if (X >= 10 && X <= 13 && Y == 34) begin oled_data = 16'hcdd1; end
    else if (X == 15 && Y == 34) begin oled_data = 16'hbd91; end
    else if (X == 16 && Y == 34) begin oled_data = 16'h840f; end
    else if (X >= 17 && X <= 32 && Y == 34) begin oled_data = 16'hcdd1; end
    else if (X == 34 && Y == 34) begin oled_data = 16'hbd91; end
    else if (X == 35 && Y == 34) begin oled_data = 16'h9cb1; end
    else if (X == 42 && Y == 34) begin oled_data = 16'hbd91; end
    else if (X == 45 && Y == 34) begin oled_data = 16'hcdd1; end
    else if (X == 46 && Y == 34) begin oled_data = 16'hbd72; end
    else if (X == 47 && Y == 34) begin oled_data = 16'h8c71; end
    else if (X == 48 && Y == 34) begin oled_data = 16'h840f; end
    else if (X == 49 && Y == 34) begin oled_data = 16'had31; end
    else if (X == 50 && Y == 34) begin oled_data = 16'hbd91; end
    else if (X >= 51 && X <= 59 && Y == 34) begin oled_data = 16'hcdd1; end
    else if (X == 60 && Y == 34) begin oled_data = 16'h8c71; end
    else if (X >= 61 && X <= 65 && Y == 34) begin oled_data = 16'hcdd1; end
    else if (X == 69 && Y == 34) begin oled_data = 16'hbd91; end
    else if (X == 71 && Y == 34) begin oled_data = 16'hcdd1; end
    else if (X == 77 && Y == 34) begin oled_data = 16'hbd91; end
    else if (X == 78 && Y == 34) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 34) begin oled_data = 16'h840f; end
    else if (X >= 80 && X <= 82 && Y == 34) begin oled_data = 16'hcdd1; end
    else if (X == 86 && Y == 34) begin oled_data = 16'hbd91; end
    else if (X == 87 && Y == 34) begin oled_data = 16'h840f; end
    else if (X == 90 && Y == 34) begin oled_data = 16'h63e9; end
    else if (X == 91 && Y == 34) begin oled_data = 16'h53c7; end
    else if (X >= 92 && X <= 93 && Y == 34) begin oled_data = 16'h5c27; end
    else if (X == 94 && Y == 34) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 34) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 35) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 35) begin oled_data = 16'h64a9; end
    else if (X == 2 && Y == 35) begin oled_data = 16'h64a9; end
    else if (X == 3 && Y == 35) begin oled_data = 16'h6468; end
    else if (X == 4 && Y == 35) begin oled_data = 16'h6468; end
    else if (X == 5 && Y == 35) begin oled_data = 16'h53c7; end
    else if (X == 6 && Y == 35) begin oled_data = 16'h740a; end
    else if (X == 7 && Y == 35) begin oled_data = 16'hcdd1; end
    else if (X == 8 && Y == 35) begin oled_data = 16'h840f; end
    else if (X >= 9 && X <= 15 && Y == 35) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 35) begin oled_data = 16'h840f; end
    else if (X == 26 && Y == 35) begin oled_data = 16'hcdd1; end
    else if (X == 34 && Y == 35) begin oled_data = 16'had31; end
    else if (X == 35 && Y == 35) begin oled_data = 16'had31; end
    else if (X == 45 && Y == 35) begin oled_data = 16'had31; end
    else if (X == 46 && Y == 35) begin oled_data = 16'h8c71; end
    else if (X == 48 && Y == 35) begin oled_data = 16'hcdd1; end
    else if (X == 49 && Y == 35) begin oled_data = 16'h8c71; end
    else if (X == 50 && Y == 35) begin oled_data = 16'had31; end
    else if (X >= 53 && X <= 59 && Y == 35) begin oled_data = 16'hcdd1; end
    else if (X == 60 && Y == 35) begin oled_data = 16'ha4f0; end
    else if (X == 61 && Y == 35) begin oled_data = 16'had31; end
    else if (X >= 69 && X <= 76 && Y == 35) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 35) begin oled_data = 16'h840f; end
    else if (X >= 80 && X <= 82 && Y == 35) begin oled_data = 16'hcdd1; end
    else if (X == 87 && Y == 35) begin oled_data = 16'h840f; end
    else if (X == 90 && Y == 35) begin oled_data = 16'h5b88; end
    else if (X == 91 && Y == 35) begin oled_data = 16'h53c7; end
    else if (X == 92 && Y == 35) begin oled_data = 16'h6468; end
    else if (X == 93 && Y == 35) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 35) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 35) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 36) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 36) begin oled_data = 16'h64a9; end
    else if (X >= 2 && X <= 4 && Y == 36) begin oled_data = 16'h5c27; end
    else if (X == 5 && Y == 36) begin oled_data = 16'h4346; end
    else if (X == 6 && Y == 36) begin oled_data = 16'ha4ee; end
    else if (X == 7 && Y == 36) begin oled_data = 16'hbd91; end
    else if (X == 8 && Y == 36) begin oled_data = 16'h840f; end
    else if (X == 9 && Y == 36) begin oled_data = 16'hcdd1; end
    else if (X == 10 && Y == 36) begin oled_data = 16'hbd91; end
    else if (X == 14 && Y == 36) begin oled_data = 16'hcdd1; end
    else if (X == 15 && Y == 36) begin oled_data = 16'hbd91; end
    else if (X == 16 && Y == 36) begin oled_data = 16'h840f; end
    else if (X >= 17 && X <= 32 && Y == 36) begin oled_data = 16'hcdd1; end
    else if (X == 34 && Y == 36) begin oled_data = 16'ha4f0; end
    else if (X == 35 && Y == 36) begin oled_data = 16'had31; end
    else if (X == 37 && Y == 36) begin oled_data = 16'hbd91; end
    else if (X == 42 && Y == 36) begin oled_data = 16'hcdd1; end
    else if (X == 45 && Y == 36) begin oled_data = 16'h8c71; end
    else if (X == 50 && Y == 36) begin oled_data = 16'h840f; end
    else if (X >= 51 && X <= 59 && Y == 36) begin oled_data = 16'hcdd1; end
    else if (X == 60 && Y == 36) begin oled_data = 16'ha4f0; end
    else if (X == 61 && Y == 36) begin oled_data = 16'ha4f0; end
    else if (X >= 65 && X <= 75 && Y == 36) begin oled_data = 16'hcdd1; end
    else if (X == 77 && Y == 36) begin oled_data = 16'hb550; end
    else if (X == 78 && Y == 36) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 36) begin oled_data = 16'h840f; end
    else if (X >= 80 && X <= 81 && Y == 36) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 36) begin oled_data = 16'hbd91; end
    else if (X == 87 && Y == 36) begin oled_data = 16'h840f; end
    else if (X >= 88 && X <= 89 && Y == 36) begin oled_data = 16'hcdd1; end
    else if (X == 90 && Y == 36) begin oled_data = 16'h4346; end
    else if (X == 91 && Y == 36) begin oled_data = 16'h53c7; end
    else if (X == 92 && Y == 36) begin oled_data = 16'h5c27; end
    else if (X == 93 && Y == 36) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 36) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 36) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 37) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 37) begin oled_data = 16'h6468; end
    else if (X == 2 && Y == 37) begin oled_data = 16'h6468; end
    else if (X == 3 && Y == 37) begin oled_data = 16'h6468; end
    else if (X == 4 && Y == 37) begin oled_data = 16'h6468; end
    else if (X == 5 && Y == 37) begin oled_data = 16'h4346; end
    else if (X == 6 && Y == 37) begin oled_data = 16'hbd91; end
    else if (X == 7 && Y == 37) begin oled_data = 16'hcdd1; end
    else if (X == 8 && Y == 37) begin oled_data = 16'h840f; end
    else if (X >= 9 && X <= 15 && Y == 37) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 37) begin oled_data = 16'h840f; end
    else if (X >= 24 && X <= 29 && Y == 37) begin oled_data = 16'hcdd1; end
    else if (X == 34 && Y == 37) begin oled_data = 16'ha4f0; end
    else if (X == 35 && Y == 37) begin oled_data = 16'hbd72; end
    else if (X == 42 && Y == 37) begin oled_data = 16'hcdd1; end
    else if (X == 45 && Y == 37) begin oled_data = 16'h8c71; end
    else if (X == 50 && Y == 37) begin oled_data = 16'h8c71; end
    else if (X >= 51 && X <= 59 && Y == 37) begin oled_data = 16'hcdd1; end
    else if (X == 60 && Y == 37) begin oled_data = 16'ha4f0; end
    else if (X == 61 && Y == 37) begin oled_data = 16'ha4f0; end
    else if (X >= 66 && X <= 67 && Y == 37) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 37) begin oled_data = 16'h840f; end
    else if (X >= 80 && X <= 85 && Y == 37) begin oled_data = 16'hcdd1; end
    else if (X == 87 && Y == 37) begin oled_data = 16'h840f; end
    else if (X == 89 && Y == 37) begin oled_data = 16'ha4ee; end
    else if (X == 90 && Y == 37) begin oled_data = 16'h4346; end
    else if (X == 91 && Y == 37) begin oled_data = 16'h5c27; end
    else if (X == 92 && Y == 37) begin oled_data = 16'h6468; end
    else if (X == 93 && Y == 37) begin oled_data = 16'h64a9; end
    else if (X == 94 && Y == 37) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 37) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 38) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 38) begin oled_data = 16'h64a9; end
    else if (X == 2 && Y == 38) begin oled_data = 16'h6468; end
    else if (X == 3 && Y == 38) begin oled_data = 16'h6468; end
    else if (X == 4 && Y == 38) begin oled_data = 16'h740a; end
    else if (X == 5 && Y == 38) begin oled_data = 16'ha4f0; end
    else if (X == 8 && Y == 38) begin oled_data = 16'h840f; end
    else if (X >= 9 && X <= 15 && Y == 38) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 38) begin oled_data = 16'h8c71; end
    else if (X >= 18 && X <= 29 && Y == 38) begin oled_data = 16'hcdd1; end
    else if (X == 34 && Y == 38) begin oled_data = 16'had31; end
    else if (X == 35 && Y == 38) begin oled_data = 16'had31; end
    else if (X == 40 && Y == 38) begin oled_data = 16'hcdd1; end
    else if (X == 45 && Y == 38) begin oled_data = 16'hbd72; end
    else if (X == 46 && Y == 38) begin oled_data = 16'h8c71; end
    else if (X == 47 && Y == 38) begin oled_data = 16'hbd72; end
    else if (X == 48 && Y == 38) begin oled_data = 16'had31; end
    else if (X == 49 && Y == 38) begin oled_data = 16'h8c71; end
    else if (X == 50 && Y == 38) begin oled_data = 16'hbd91; end
    else if (X >= 52 && X <= 59 && Y == 38) begin oled_data = 16'hcdd1; end
    else if (X == 60 && Y == 38) begin oled_data = 16'ha4f0; end
    else if (X == 61 && Y == 38) begin oled_data = 16'had31; end
    else if (X >= 66 && X <= 68 && Y == 38) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 38) begin oled_data = 16'h840f; end
    else if (X >= 80 && X <= 86 && Y == 38) begin oled_data = 16'hcdd1; end
    else if (X == 87 && Y == 38) begin oled_data = 16'h73af; end
    else if (X == 88 && Y == 38) begin oled_data = 16'hcdd1; end
    else if (X == 89 && Y == 38) begin oled_data = 16'h848c; end
    else if (X == 90 && Y == 38) begin oled_data = 16'h4346; end
    else if (X == 91 && Y == 38) begin oled_data = 16'h53c7; end
    else if (X == 92 && Y == 38) begin oled_data = 16'h5c27; end
    else if (X == 93 && Y == 38) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 38) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 38) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 39) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 39) begin oled_data = 16'h64a9; end
    else if (X == 2 && Y == 39) begin oled_data = 16'h6468; end
    else if (X == 3 && Y == 39) begin oled_data = 16'h64a9; end
    else if (X == 4 && Y == 39) begin oled_data = 16'h6468; end
    else if (X == 5 && Y == 39) begin oled_data = 16'h848c; end
    else if (X == 8 && Y == 39) begin oled_data = 16'h8c71; end
    else if (X == 9 && Y == 39) begin oled_data = 16'hb550; end
    else if (X >= 13 && X <= 14 && Y == 39) begin oled_data = 16'hcdd1; end
    else if (X == 15 && Y == 39) begin oled_data = 16'hbd91; end
    else if (X == 16 && Y == 39) begin oled_data = 16'h8c71; end
    else if (X >= 22 && X <= 33 && Y == 39) begin oled_data = 16'hcdd1; end
    else if (X == 34 && Y == 39) begin oled_data = 16'hbd91; end
    else if (X == 35 && Y == 39) begin oled_data = 16'h8c71; end
    else if (X == 46 && Y == 39) begin oled_data = 16'hc5d3; end
    else if (X == 47 && Y == 39) begin oled_data = 16'h94b2; end
    else if (X == 48 && Y == 39) begin oled_data = 16'h8c71; end
    else if (X == 49 && Y == 39) begin oled_data = 16'hbd91; end
    else if (X == 50 && Y == 39) begin oled_data = 16'hbd91; end
    else if (X >= 51 && X <= 56 && Y == 39) begin oled_data = 16'hcdd1; end
    else if (X == 58 && Y == 39) begin oled_data = 16'hbd91; end
    else if (X == 59 && Y == 39) begin oled_data = 16'hcdd1; end
    else if (X == 60 && Y == 39) begin oled_data = 16'h8c71; end
    else if (X == 61 && Y == 39) begin oled_data = 16'hc5b2; end
    else if (X >= 65 && X <= 78 && Y == 39) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 39) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 39) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 39) begin oled_data = 16'hb550; end
    else if (X >= 83 && X <= 85 && Y == 39) begin oled_data = 16'hcdd1; end
    else if (X == 86 && Y == 39) begin oled_data = 16'had0f; end
    else if (X == 87 && Y == 39) begin oled_data = 16'h8c71; end
    else if (X == 88 && Y == 39) begin oled_data = 16'hcdd1; end
    else if (X == 89 && Y == 39) begin oled_data = 16'h5bc8; end
    else if (X == 90 && Y == 39) begin oled_data = 16'h4346; end
    else if (X == 91 && Y == 39) begin oled_data = 16'h53c7; end
    else if (X >= 92 && X <= 93 && Y == 39) begin oled_data = 16'h5c27; end
    else if (X == 94 && Y == 39) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 39) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 40) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 40) begin oled_data = 16'h64a9; end
    else if (X == 2 && Y == 40) begin oled_data = 16'h64a9; end
    else if (X == 3 && Y == 40) begin oled_data = 16'h64a9; end
    else if (X == 4 && Y == 40) begin oled_data = 16'h64a9; end
    else if (X == 5 && Y == 40) begin oled_data = 16'h53c7; end
    else if (X == 6 && Y == 40) begin oled_data = 16'h7c4b; end
    else if (X == 7 && Y == 40) begin oled_data = 16'had0f; end
    else if (X == 8 && Y == 40) begin oled_data = 16'hbd91; end
    else if (X == 9 && Y == 40) begin oled_data = 16'h840f; end
    else if (X >= 10 && X <= 13 && Y == 40) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 40) begin oled_data = 16'h8c71; end
    else if (X == 35 && Y == 40) begin oled_data = 16'h840f; end
    else if (X == 38 && Y == 40) begin oled_data = 16'hde75; end
    else if (X == 39 && Y == 40) begin oled_data = 16'hde75; end
    else if (X == 40 && Y == 40) begin oled_data = 16'hde75; end
    else if (X == 41 && Y == 40) begin oled_data = 16'hde75; end
    else if (X == 42 && Y == 40) begin oled_data = 16'hde75; end
    else if (X == 47 && Y == 40) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 40) begin oled_data = 16'had31; end
    else if (X >= 51 && X <= 56 && Y == 40) begin oled_data = 16'hcdd1; end
    else if (X == 60 && Y == 40) begin oled_data = 16'h840f; end
    else if (X >= 66 && X <= 75 && Y == 40) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 40) begin oled_data = 16'h840f; end
    else if (X >= 80 && X <= 85 && Y == 40) begin oled_data = 16'hcdd1; end
    else if (X == 86 && Y == 40) begin oled_data = 16'h840f; end
    else if (X == 87 && Y == 40) begin oled_data = 16'hcdd1; end
    else if (X == 88 && Y == 40) begin oled_data = 16'ha4ee; end
    else if (X == 89 && Y == 40) begin oled_data = 16'h53c7; end
    else if (X == 90 && Y == 40) begin oled_data = 16'h4346; end
    else if (X == 91 && Y == 40) begin oled_data = 16'h53c7; end
    else if (X == 92 && Y == 40) begin oled_data = 16'h5c27; end
    else if (X == 93 && Y == 40) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 40) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 40) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 41) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 41) begin oled_data = 16'h64a9; end
    else if (X == 2 && Y == 41) begin oled_data = 16'h6468; end
    else if (X == 3 && Y == 41) begin oled_data = 16'h64a9; end
    else if (X == 4 && Y == 41) begin oled_data = 16'h6468; end
    else if (X == 5 && Y == 41) begin oled_data = 16'h53c7; end
    else if (X == 6 && Y == 41) begin oled_data = 16'h5c27; end
    else if (X == 7 && Y == 41) begin oled_data = 16'h53c7; end
    else if (X == 8 && Y == 41) begin oled_data = 16'h740a; end
    else if (X == 9 && Y == 41) begin oled_data = 16'ha4f0; end
    else if (X == 10 && Y == 41) begin oled_data = 16'h8c71; end
    else if (X >= 11 && X <= 15 && Y == 41) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 41) begin oled_data = 16'h840f; end
    else if (X >= 17 && X <= 34 && Y == 41) begin oled_data = 16'hcdd1; end
    else if (X == 35 && Y == 41) begin oled_data = 16'h9cb1; end
    else if (X == 36 && Y == 41) begin oled_data = 16'had31; end
    else if (X == 37 && Y == 41) begin oled_data = 16'hcdd1; end
    else if (X == 42 && Y == 41) begin oled_data = 16'hc5b2; end
    else if (X == 47 && Y == 41) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 41) begin oled_data = 16'ha4f0; end
    else if (X >= 49 && X <= 58 && Y == 41) begin oled_data = 16'hcdd1; end
    else if (X == 59 && Y == 41) begin oled_data = 16'ha4f0; end
    else if (X == 60 && Y == 41) begin oled_data = 16'h9cb1; end
    else if (X >= 61 && X <= 65 && Y == 41) begin oled_data = 16'hcdd1; end
    else if (X == 66 && Y == 41) begin oled_data = 16'hbd91; end
    else if (X >= 67 && X <= 75 && Y == 41) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 41) begin oled_data = 16'h840f; end
    else if (X >= 80 && X <= 83 && Y == 41) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 41) begin oled_data = 16'h840f; end
    else if (X == 86 && Y == 41) begin oled_data = 16'ha4f0; end
    else if (X == 87 && Y == 41) begin oled_data = 16'hb550; end
    else if (X == 88 && Y == 41) begin oled_data = 16'h5bc8; end
    else if (X == 89 && Y == 41) begin oled_data = 16'h53c7; end
    else if (X == 90 && Y == 41) begin oled_data = 16'h4346; end
    else if (X == 91 && Y == 41) begin oled_data = 16'h53c7; end
    else if (X >= 92 && X <= 93 && Y == 41) begin oled_data = 16'h5c27; end
    else if (X == 94 && Y == 41) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 41) begin oled_data = 16'h9551; end
    else if (X == 0 && Y == 42) begin oled_data = 16'hadd4; end
    else if (X == 1 && Y == 42) begin oled_data = 16'h6468; end
    else if (X == 2 && Y == 42) begin oled_data = 16'h64a9; end
    else if (X == 3 && Y == 42) begin oled_data = 16'h7509; end
    else if (X == 4 && Y == 42) begin oled_data = 16'h64a9; end
    else if (X == 5 && Y == 42) begin oled_data = 16'h5c27; end
    else if (X == 6 && Y == 42) begin oled_data = 16'h6468; end
    else if (X == 7 && Y == 42) begin oled_data = 16'h5c27; end
    else if (X == 8 && Y == 42) begin oled_data = 16'h53c7; end
    else if (X == 9 && Y == 42) begin oled_data = 16'h9cad; end
    else if (X == 10 && Y == 42) begin oled_data = 16'h9c8e; end
    else if (X == 11 && Y == 42) begin oled_data = 16'h840f; end
    else if (X >= 12 && X <= 15 && Y == 42) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 42) begin oled_data = 16'h8c71; end
    else if (X >= 17 && X <= 18 && Y == 42) begin oled_data = 16'hcdd1; end
    else if (X == 36 && Y == 42) begin oled_data = 16'h8c71; end
    else if (X == 40 && Y == 42) begin oled_data = 16'hde75; end
    else if (X == 41 && Y == 42) begin oled_data = 16'hde75; end
    else if (X == 42 && Y == 42) begin oled_data = 16'hde75; end
    else if (X == 43 && Y == 42) begin oled_data = 16'hde75; end
    else if (X == 44 && Y == 42) begin oled_data = 16'hde75; end
    else if (X == 47 && Y == 42) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 42) begin oled_data = 16'had31; end
    else if (X >= 49 && X <= 58 && Y == 42) begin oled_data = 16'hcdd1; end
    else if (X == 59 && Y == 42) begin oled_data = 16'h8c71; end
    else if (X == 72 && Y == 42) begin oled_data = 16'hde75; end
    else if (X == 79 && Y == 42) begin oled_data = 16'h840f; end
    else if (X == 83 && Y == 42) begin oled_data = 16'hbd91; end
    else if (X == 84 && Y == 42) begin oled_data = 16'h840f; end
    else if (X == 85 && Y == 42) begin oled_data = 16'ha4f0; end
    else if (X == 87 && Y == 42) begin oled_data = 16'h848c; end
    else if (X == 88 && Y == 42) begin oled_data = 16'h6468; end
    else if (X == 89 && Y == 42) begin oled_data = 16'h5c27; end
    else if (X == 90 && Y == 42) begin oled_data = 16'h4346; end
    else if (X == 91 && Y == 42) begin oled_data = 16'h53c7; end
    else if (X == 92 && Y == 42) begin oled_data = 16'h6468; end
    else if (X == 93 && Y == 42) begin oled_data = 16'h64a9; end
    else if (X == 94 && Y == 42) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 42) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 43) begin oled_data = 16'hadd4; end
    else if (X == 1 && Y == 43) begin oled_data = 16'h64a9; end
    else if (X == 2 && Y == 43) begin oled_data = 16'h64a9; end
    else if (X == 3 && Y == 43) begin oled_data = 16'h7509; end
    else if (X == 4 && Y == 43) begin oled_data = 16'h7509; end
    else if (X == 5 && Y == 43) begin oled_data = 16'h5c27; end
    else if (X == 6 && Y == 43) begin oled_data = 16'h6468; end
    else if (X == 7 && Y == 43) begin oled_data = 16'h5c27; end
    else if (X == 8 && Y == 43) begin oled_data = 16'h53c7; end
    else if (X == 9 && Y == 43) begin oled_data = 16'h740a; end
    else if (X == 10 && Y == 43) begin oled_data = 16'hcdd1; end
    else if (X == 11 && Y == 43) begin oled_data = 16'hbd91; end
    else if (X == 12 && Y == 43) begin oled_data = 16'h840f; end
    else if (X == 13 && Y == 43) begin oled_data = 16'h840f; end
    else if (X == 14 && Y == 43) begin oled_data = 16'ha4f0; end
    else if (X == 15 && Y == 43) begin oled_data = 16'ha4f0; end
    else if (X == 16 && Y == 43) begin oled_data = 16'h840f; end
    else if (X == 17 && Y == 43) begin oled_data = 16'hcdd1; end
    else if (X == 29 && Y == 43) begin oled_data = 16'hde75; end
    else if (X == 36 && Y == 43) begin oled_data = 16'had31; end
    else if (X == 37 && Y == 43) begin oled_data = 16'had31; end
    else if (X == 42 && Y == 43) begin oled_data = 16'hde75; end
    else if (X == 43 && Y == 43) begin oled_data = 16'hde75; end
    else if (X == 44 && Y == 43) begin oled_data = 16'hde75; end
    else if (X == 47 && Y == 43) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 43) begin oled_data = 16'had31; end
    else if (X >= 49 && X <= 55 && Y == 43) begin oled_data = 16'hcdd1; end
    else if (X == 58 && Y == 43) begin oled_data = 16'ha4f0; end
    else if (X == 59 && Y == 43) begin oled_data = 16'had31; end
    else if (X == 65 && Y == 43) begin oled_data = 16'hde75; end
    else if (X == 69 && Y == 43) begin oled_data = 16'hde75; end
    else if (X == 75 && Y == 43) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 43) begin oled_data = 16'h8c71; end
    else if (X == 80 && Y == 43) begin oled_data = 16'ha4f0; end
    else if (X == 81 && Y == 43) begin oled_data = 16'ha4f0; end
    else if (X == 82 && Y == 43) begin oled_data = 16'h840f; end
    else if (X == 83 && Y == 43) begin oled_data = 16'h8c71; end
    else if (X == 84 && Y == 43) begin oled_data = 16'hcdd1; end
    else if (X == 86 && Y == 43) begin oled_data = 16'had31; end
    else if (X == 87 && Y == 43) begin oled_data = 16'h5c27; end
    else if (X == 88 && Y == 43) begin oled_data = 16'h6468; end
    else if (X == 89 && Y == 43) begin oled_data = 16'h5c27; end
    else if (X == 90 && Y == 43) begin oled_data = 16'h4346; end
    else if (X >= 91 && X <= 92 && Y == 43) begin oled_data = 16'h5c27; end
    else if (X == 93 && Y == 43) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 43) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 43) begin oled_data = 16'hadd4; end
    else if (X == 0 && Y == 44) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 44) begin oled_data = 16'h6468; end
    else if (X == 2 && Y == 44) begin oled_data = 16'h6468; end
    else if (X == 3 && Y == 44) begin oled_data = 16'h6468; end
    else if (X == 4 && Y == 44) begin oled_data = 16'h64a9; end
    else if (X == 5 && Y == 44) begin oled_data = 16'h53c7; end
    else if (X == 6 && Y == 44) begin oled_data = 16'h6468; end
    else if (X == 7 && Y == 44) begin oled_data = 16'h5c27; end
    else if (X == 8 && Y == 44) begin oled_data = 16'h53c7; end
    else if (X == 9 && Y == 44) begin oled_data = 16'h53c7; end
    else if (X == 10 && Y == 44) begin oled_data = 16'ha4ee; end
    else if (X == 11 && Y == 44) begin oled_data = 16'hcdd1; end
    else if (X == 13 && Y == 44) begin oled_data = 16'hb550; end
    else if (X == 14 && Y == 44) begin oled_data = 16'had0f; end
    else if (X == 15 && Y == 44) begin oled_data = 16'h8c71; end
    else if (X == 16 && Y == 44) begin oled_data = 16'h840f; end
    else if (X >= 17 && X <= 29 && Y == 44) begin oled_data = 16'hcdd1; end
    else if (X == 37 && Y == 44) begin oled_data = 16'h8c71; end
    else if (X == 38 && Y == 44) begin oled_data = 16'had31; end
    else if (X == 39 && Y == 44) begin oled_data = 16'hcdd1; end
    else if (X == 42 && Y == 44) begin oled_data = 16'hc5d3; end
    else if (X == 43 && Y == 44) begin oled_data = 16'hde75; end
    else if (X == 44 && Y == 44) begin oled_data = 16'hde75; end
    else if (X == 45 && Y == 44) begin oled_data = 16'hc5b2; end
    else if (X == 47 && Y == 44) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 44) begin oled_data = 16'ha4f0; end
    else if (X == 49 && Y == 44) begin oled_data = 16'hcdd1; end
    else if (X == 50 && Y == 44) begin oled_data = 16'hb550; end
    else if (X >= 51 && X <= 56 && Y == 44) begin oled_data = 16'hcdd1; end
    else if (X == 57 && Y == 44) begin oled_data = 16'ha4f0; end
    else if (X == 58 && Y == 44) begin oled_data = 16'h9cb1; end
    else if (X >= 60 && X <= 77 && Y == 44) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 44) begin oled_data = 16'h8c71; end
    else if (X == 80 && Y == 44) begin oled_data = 16'ha4f0; end
    else if (X == 81 && Y == 44) begin oled_data = 16'had31; end
    else if (X == 82 && Y == 44) begin oled_data = 16'hbd91; end
    else if (X == 83 && Y == 44) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 44) begin oled_data = 16'h9cad; end
    else if (X >= 86 && X <= 89 && Y == 44) begin oled_data = 16'h5c27; end
    else if (X == 90 && Y == 44) begin oled_data = 16'h4346; end
    else if (X == 91 && Y == 44) begin oled_data = 16'h53c7; end
    else if (X == 92 && Y == 44) begin oled_data = 16'h5c27; end
    else if (X == 93 && Y == 44) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 44) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 44) begin oled_data = 16'hb5b6; end
    else if (X == 0 && Y == 45) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 45) begin oled_data = 16'h64a9; end
    else if (X == 2 && Y == 45) begin oled_data = 16'h64a9; end
    else if (X == 3 && Y == 45) begin oled_data = 16'h7509; end
    else if (X == 4 && Y == 45) begin oled_data = 16'h64a9; end
    else if (X == 5 && Y == 45) begin oled_data = 16'h5c27; end
    else if (X == 6 && Y == 45) begin oled_data = 16'h64a9; end
    else if (X == 7 && Y == 45) begin oled_data = 16'h64a9; end
    else if (X >= 8 && X <= 9 && Y == 45) begin oled_data = 16'h5c27; end
    else if (X == 10 && Y == 45) begin oled_data = 16'h53c7; end
    else if (X >= 11 && X <= 15 && Y == 45) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 45) begin oled_data = 16'h840f; end
    else if (X >= 17 && X <= 18 && Y == 45) begin oled_data = 16'hcdd1; end
    else if (X == 31 && Y == 45) begin oled_data = 16'hde75; end
    else if (X == 38 && Y == 45) begin oled_data = 16'h8c71; end
    else if (X == 39 && Y == 45) begin oled_data = 16'had31; end
    else if (X == 41 && Y == 45) begin oled_data = 16'hde75; end
    else if (X == 42 && Y == 45) begin oled_data = 16'hde75; end
    else if (X == 43 && Y == 45) begin oled_data = 16'hde75; end
    else if (X == 44 && Y == 45) begin oled_data = 16'hde75; end
    else if (X == 45 && Y == 45) begin oled_data = 16'hde75; end
    else if (X == 47 && Y == 45) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 45) begin oled_data = 16'had31; end
    else if (X >= 49 && X <= 55 && Y == 45) begin oled_data = 16'hcdd1; end
    else if (X == 56 && Y == 45) begin oled_data = 16'ha4f0; end
    else if (X == 57 && Y == 45) begin oled_data = 16'h8c71; end
    else if (X == 65 && Y == 45) begin oled_data = 16'hde75; end
    else if (X >= 69 && X <= 77 && Y == 45) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 45) begin oled_data = 16'h8c71; end
    else if (X >= 80 && X <= 82 && Y == 45) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 45) begin oled_data = 16'h740a; end
    else if (X == 86 && Y == 45) begin oled_data = 16'h6468; end
    else if (X == 87 && Y == 45) begin oled_data = 16'h6468; end
    else if (X == 88 && Y == 45) begin oled_data = 16'h6468; end
    else if (X == 89 && Y == 45) begin oled_data = 16'h5c27; end
    else if (X == 90 && Y == 45) begin oled_data = 16'h4346; end
    else if (X == 91 && Y == 45) begin oled_data = 16'h5c27; end
    else if (X == 92 && Y == 45) begin oled_data = 16'h64a9; end
    else if (X == 93 && Y == 45) begin oled_data = 16'h64a9; end
    else if (X == 94 && Y == 45) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 45) begin oled_data = 16'hb5b6; end
    else if (X == 0 && Y == 46) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 46) begin oled_data = 16'h64a9; end
    else if (X == 2 && Y == 46) begin oled_data = 16'h64a9; end
    else if (X == 3 && Y == 46) begin oled_data = 16'h64a9; end
    else if (X == 4 && Y == 46) begin oled_data = 16'h6468; end
    else if (X == 5 && Y == 46) begin oled_data = 16'h5b88; end
    else if (X >= 6 && X <= 7 && Y == 46) begin oled_data = 16'h5c27; end
    else if (X == 8 && Y == 46) begin oled_data = 16'h53c7; end
    else if (X == 9 && Y == 46) begin oled_data = 16'h53c7; end
    else if (X == 10 && Y == 46) begin oled_data = 16'h4b07; end
    else if (X == 11 && Y == 46) begin oled_data = 16'had0f; end
    else if (X == 12 && Y == 46) begin oled_data = 16'hb550; end
    else if (X == 13 && Y == 46) begin oled_data = 16'ha4f0; end
    else if (X == 15 && Y == 46) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 46) begin oled_data = 16'h840f; end
    else if (X == 17 && Y == 46) begin oled_data = 16'hcdd1; end
    else if (X == 18 && Y == 46) begin oled_data = 16'hbd91; end
    else if (X >= 22 && X <= 28 && Y == 46) begin oled_data = 16'hcdd1; end
    else if (X == 39 && Y == 46) begin oled_data = 16'h9cb1; end
    else if (X == 40 && Y == 46) begin oled_data = 16'h9cb1; end
    else if (X == 41 && Y == 46) begin oled_data = 16'hcdd1; end
    else if (X == 45 && Y == 46) begin oled_data = 16'hc5d3; end
    else if (X == 47 && Y == 46) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 46) begin oled_data = 16'had31; end
    else if (X >= 50 && X <= 54 && Y == 46) begin oled_data = 16'hcdd1; end
    else if (X == 55 && Y == 46) begin oled_data = 16'h8c71; end
    else if (X == 56 && Y == 46) begin oled_data = 16'h9cb1; end
    else if (X >= 61 && X <= 78 && Y == 46) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 46) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 46) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 46) begin oled_data = 16'h9c8e; end
    else if (X == 83 && Y == 46) begin oled_data = 16'hb550; end
    else if (X == 84 && Y == 46) begin oled_data = 16'h9cad; end
    else if (X == 85 && Y == 46) begin oled_data = 16'h4346; end
    else if (X == 86 && Y == 46) begin oled_data = 16'h53c7; end
    else if (X == 87 && Y == 46) begin oled_data = 16'h53c7; end
    else if (X == 88 && Y == 46) begin oled_data = 16'h53c7; end
    else if (X == 89 && Y == 46) begin oled_data = 16'h53c7; end
    else if (X == 90 && Y == 46) begin oled_data = 16'h4b07; end
    else if (X == 91 && Y == 46) begin oled_data = 16'h5c27; end
    else if (X == 92 && Y == 46) begin oled_data = 16'h6468; end
    else if (X == 93 && Y == 46) begin oled_data = 16'h5c27; end
    else if (X == 94 && Y == 46) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 46) begin oled_data = 16'hadd4; end
    else if (X == 0 && Y == 47) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 47) begin oled_data = 16'h7509; end
    else if (X == 2 && Y == 47) begin oled_data = 16'h7509; end
    else if (X == 3 && Y == 47) begin oled_data = 16'h7509; end
    else if (X == 4 && Y == 47) begin oled_data = 16'h64a9; end
    else if (X == 5 && Y == 47) begin oled_data = 16'h6468; end
    else if (X == 6 && Y == 47) begin oled_data = 16'h64a9; end
    else if (X == 7 && Y == 47) begin oled_data = 16'h64a9; end
    else if (X == 8 && Y == 47) begin oled_data = 16'h5c27; end
    else if (X == 9 && Y == 47) begin oled_data = 16'h538c; end
    else if (X == 10 && Y == 47) begin oled_data = 16'h4b07; end
    else if (X >= 11 && X <= 13 && Y == 47) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 47) begin oled_data = 16'h8c71; end
    else if (X >= 17 && X <= 26 && Y == 47) begin oled_data = 16'hcdd1; end
    else if (X == 40 && Y == 47) begin oled_data = 16'hc5b2; end
    else if (X == 41 && Y == 47) begin oled_data = 16'h8c71; end
    else if (X == 42 && Y == 47) begin oled_data = 16'h9cb1; end
    else if (X == 47 && Y == 47) begin oled_data = 16'hb573; end
    else if (X == 48 && Y == 47) begin oled_data = 16'had31; end
    else if (X == 52 && Y == 47) begin oled_data = 16'hcdd1; end
    else if (X == 53 && Y == 47) begin oled_data = 16'h9cb1; end
    else if (X == 54 && Y == 47) begin oled_data = 16'h8c71; end
    else if (X == 55 && Y == 47) begin oled_data = 16'hc5b2; end
    else if (X == 58 && Y == 47) begin oled_data = 16'hcdd1; end
    else if (X == 72 && Y == 47) begin oled_data = 16'hde75; end
    else if (X == 79 && Y == 47) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 47) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 47) begin oled_data = 16'hb550; end
    else if (X == 84 && Y == 47) begin oled_data = 16'h9cad; end
    else if (X >= 85 && X <= 91 && Y == 47) begin oled_data = 16'h5c27; end
    else if (X == 92 && Y == 47) begin oled_data = 16'h6468; end
    else if (X == 93 && Y == 47) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 47) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 47) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 48) begin oled_data = 16'h9551; end
    else if (X == 1 && Y == 48) begin oled_data = 16'h7509; end
    else if (X == 2 && Y == 48) begin oled_data = 16'h7509; end
    else if (X == 3 && Y == 48) begin oled_data = 16'h64a9; end
    else if (X == 4 && Y == 48) begin oled_data = 16'h64a9; end
    else if (X == 5 && Y == 48) begin oled_data = 16'h64a9; end
    else if (X == 6 && Y == 48) begin oled_data = 16'h64a9; end
    else if (X == 7 && Y == 48) begin oled_data = 16'h6468; end
    else if (X == 8 && Y == 48) begin oled_data = 16'h53c7; end
    else if (X == 9 && Y == 48) begin oled_data = 16'h5b88; end
    else if (X == 10 && Y == 48) begin oled_data = 16'h4b07; end
    else if (X >= 13 && X <= 15 && Y == 48) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 48) begin oled_data = 16'h8c71; end
    else if (X >= 17 && X <= 26 && Y == 48) begin oled_data = 16'hcdd1; end
    else if (X == 30 && Y == 48) begin oled_data = 16'hde75; end
    else if (X == 33 && Y == 48) begin oled_data = 16'hde75; end
    else if (X == 36 && Y == 48) begin oled_data = 16'hde75; end
    else if (X == 42 && Y == 48) begin oled_data = 16'had31; end
    else if (X == 43 && Y == 48) begin oled_data = 16'h94b2; end
    else if (X == 44 && Y == 48) begin oled_data = 16'h8c71; end
    else if (X == 45 && Y == 48) begin oled_data = 16'h94b2; end
    else if (X == 46 && Y == 48) begin oled_data = 16'hb573; end
    else if (X == 47 && Y == 48) begin oled_data = 16'h94b2; end
    else if (X == 48 && Y == 48) begin oled_data = 16'h8c71; end
    else if (X == 49 && Y == 48) begin oled_data = 16'ha4f0; end
    else if (X == 50 && Y == 48) begin oled_data = 16'h8c71; end
    else if (X == 51 && Y == 48) begin oled_data = 16'h8c71; end
    else if (X == 52 && Y == 48) begin oled_data = 16'h94b2; end
    else if (X == 53 && Y == 48) begin oled_data = 16'hbd72; end
    else if (X >= 58 && X <= 77 && Y == 48) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 48) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 48) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 48) begin oled_data = 16'hb550; end
    else if (X == 84 && Y == 48) begin oled_data = 16'hbd91; end
    else if (X >= 85 && X <= 90 && Y == 48) begin oled_data = 16'h5c27; end
    else if (X == 91 && Y == 48) begin oled_data = 16'h6468; end
    else if (X == 92 && Y == 48) begin oled_data = 16'h6468; end
    else if (X == 93 && Y == 48) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 48) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 48) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 49) begin oled_data = 16'h9551; end
    else if (X == 1 && Y == 49) begin oled_data = 16'h6468; end
    else if (X == 2 && Y == 49) begin oled_data = 16'h6468; end
    else if (X == 3 && Y == 49) begin oled_data = 16'h64a9; end
    else if (X == 4 && Y == 49) begin oled_data = 16'h7509; end
    else if (X == 5 && Y == 49) begin oled_data = 16'h6468; end
    else if (X == 6 && Y == 49) begin oled_data = 16'h6468; end
    else if (X == 7 && Y == 49) begin oled_data = 16'h5c27; end
    else if (X == 8 && Y == 49) begin oled_data = 16'h53c7; end
    else if (X == 9 && Y == 49) begin oled_data = 16'h52ca; end
    else if (X == 10 && Y == 49) begin oled_data = 16'h4b07; end
    else if (X == 11 && Y == 49) begin oled_data = 16'hcdd1; end
    else if (X == 13 && Y == 49) begin oled_data = 16'h9c8e; end
    else if (X == 15 && Y == 49) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 49) begin oled_data = 16'h8c71; end
    else if (X >= 17 && X <= 28 && Y == 49) begin oled_data = 16'hcdd1; end
    else if (X == 30 && Y == 49) begin oled_data = 16'hc5d3; end
    else if (X == 34 && Y == 49) begin oled_data = 16'hbd91; end
    else if (X >= 35 && X <= 45 && Y == 49) begin oled_data = 16'hcdd1; end
    else if (X == 46 && Y == 49) begin oled_data = 16'hbd72; end
    else if (X == 47 && Y == 49) begin oled_data = 16'h8c71; end
    else if (X == 48 && Y == 49) begin oled_data = 16'h9cb1; end
    else if (X == 49 && Y == 49) begin oled_data = 16'hbd72; end
    else if (X >= 50 && X <= 60 && Y == 49) begin oled_data = 16'hcdd1; end
    else if (X == 61 && Y == 49) begin oled_data = 16'hb550; end
    else if (X >= 62 && X <= 76 && Y == 49) begin oled_data = 16'hcdd1; end
    else if (X == 77 && Y == 49) begin oled_data = 16'hbd91; end
    else if (X == 78 && Y == 49) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 49) begin oled_data = 16'h840f; end
    else if (X == 82 && Y == 49) begin oled_data = 16'hb550; end
    else if (X == 84 && Y == 49) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 49) begin oled_data = 16'h53c7; end
    else if (X >= 86 && X <= 88 && Y == 49) begin oled_data = 16'h5c27; end
    else if (X == 89 && Y == 49) begin oled_data = 16'h6468; end
    else if (X == 90 && Y == 49) begin oled_data = 16'h5c27; end
    else if (X == 91 && Y == 49) begin oled_data = 16'h6468; end
    else if (X == 92 && Y == 49) begin oled_data = 16'h64a9; end
    else if (X == 93 && Y == 49) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 49) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 49) begin oled_data = 16'h9551; end
    else if (X == 0 && Y == 50) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 50) begin oled_data = 16'h6468; end
    else if (X == 2 && Y == 50) begin oled_data = 16'h6468; end
    else if (X == 3 && Y == 50) begin oled_data = 16'h64a9; end
    else if (X == 4 && Y == 50) begin oled_data = 16'h7509; end
    else if (X == 5 && Y == 50) begin oled_data = 16'h6468; end
    else if (X == 6 && Y == 50) begin oled_data = 16'h64a9; end
    else if (X == 7 && Y == 50) begin oled_data = 16'h5c27; end
    else if (X == 8 && Y == 50) begin oled_data = 16'h53c7; end
    else if (X == 9 && Y == 50) begin oled_data = 16'h5c27; end
    else if (X == 10 && Y == 50) begin oled_data = 16'h4346; end
    else if (X == 11 && Y == 50) begin oled_data = 16'hcdd1; end
    else if (X == 13 && Y == 50) begin oled_data = 16'hb550; end
    else if (X == 15 && Y == 50) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 50) begin oled_data = 16'h8c71; end
    else if (X >= 17 && X <= 34 && Y == 50) begin oled_data = 16'hcdd1; end
    else if (X == 47 && Y == 50) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 50) begin oled_data = 16'had31; end
    else if (X >= 74 && X <= 78 && Y == 50) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 50) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 50) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 50) begin oled_data = 16'hb550; end
    else if (X == 85 && Y == 50) begin oled_data = 16'h7c4b; end
    else if (X >= 86 && X <= 88 && Y == 50) begin oled_data = 16'h5c27; end
    else if (X == 89 && Y == 50) begin oled_data = 16'h6468; end
    else if (X == 90 && Y == 50) begin oled_data = 16'h64a9; end
    else if (X == 91 && Y == 50) begin oled_data = 16'h7509; end
    else if (X == 92 && Y == 50) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 50) begin oled_data = 16'h7509; end
    else if (X == 94 && Y == 50) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 50) begin oled_data = 16'h9551; end
    else if (X == 0 && Y == 51) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 51) begin oled_data = 16'h53c7; end
    else if (X >= 2 && X <= 3 && Y == 51) begin oled_data = 16'h5c27; end
    else if (X == 4 && Y == 51) begin oled_data = 16'h6468; end
    else if (X == 5 && Y == 51) begin oled_data = 16'h5c27; end
    else if (X == 6 && Y == 51) begin oled_data = 16'h6468; end
    else if (X == 7 && Y == 51) begin oled_data = 16'h5c27; end
    else if (X == 8 && Y == 51) begin oled_data = 16'h53c7; end
    else if (X == 9 && Y == 51) begin oled_data = 16'h5c27; end
    else if (X == 10 && Y == 51) begin oled_data = 16'h4346; end
    else if (X == 11 && Y == 51) begin oled_data = 16'hbd91; end
    else if (X == 13 && Y == 51) begin oled_data = 16'had0f; end
    else if (X == 15 && Y == 51) begin oled_data = 16'hbd91; end
    else if (X == 16 && Y == 51) begin oled_data = 16'h840f; end
    else if (X == 17 && Y == 51) begin oled_data = 16'hcdd1; end
    else if (X == 18 && Y == 51) begin oled_data = 16'hbd91; end
    else if (X >= 24 && X <= 46 && Y == 51) begin oled_data = 16'hcdd1; end
    else if (X == 47 && Y == 51) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 51) begin oled_data = 16'had31; end
    else if (X == 50 && Y == 51) begin oled_data = 16'hbd91; end
    else if (X >= 52 && X <= 69 && Y == 51) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 51) begin oled_data = 16'h840f; end
    else if (X >= 80 && X <= 81 && Y == 51) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 51) begin oled_data = 16'had0f; end
    else if (X == 85 && Y == 51) begin oled_data = 16'hb550; end
    else if (X == 86 && Y == 51) begin oled_data = 16'h7c4b; end
    else if (X == 87 && Y == 51) begin oled_data = 16'h53c7; end
    else if (X == 88 && Y == 51) begin oled_data = 16'h5c27; end
    else if (X == 89 && Y == 51) begin oled_data = 16'h6468; end
    else if (X == 90 && Y == 51) begin oled_data = 16'h6468; end
    else if (X == 91 && Y == 51) begin oled_data = 16'h7509; end
    else if (X == 92 && Y == 51) begin oled_data = 16'h7509; end
    else if (X == 93 && Y == 51) begin oled_data = 16'h64a9; end
    else if (X == 94 && Y == 51) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 51) begin oled_data = 16'h9551; end
    else if (X == 0 && Y == 52) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 52) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 52) begin oled_data = 16'h6468; end
    else if (X == 3 && Y == 52) begin oled_data = 16'h64a9; end
    else if (X == 4 && Y == 52) begin oled_data = 16'h64a9; end
    else if (X == 5 && Y == 52) begin oled_data = 16'h5c27; end
    else if (X == 6 && Y == 52) begin oled_data = 16'h64a9; end
    else if (X == 7 && Y == 52) begin oled_data = 16'h6468; end
    else if (X >= 8 && X <= 9 && Y == 52) begin oled_data = 16'h5c27; end
    else if (X == 10 && Y == 52) begin oled_data = 16'h53c7; end
    else if (X == 11 && Y == 52) begin oled_data = 16'hcdd1; end
    else if (X == 13 && Y == 52) begin oled_data = 16'hb550; end
    else if (X == 15 && Y == 52) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 52) begin oled_data = 16'h8c71; end
    else if (X >= 17 && X <= 23 && Y == 52) begin oled_data = 16'hcdd1; end
    else if (X == 47 && Y == 52) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 52) begin oled_data = 16'had31; end
    else if (X >= 61 && X <= 67 && Y == 52) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 52) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 52) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 52) begin oled_data = 16'hb550; end
    else if (X == 87 && Y == 52) begin oled_data = 16'h848c; end
    else if (X == 88 && Y == 52) begin oled_data = 16'h5c27; end
    else if (X == 89 && Y == 52) begin oled_data = 16'h64a9; end
    else if (X == 90 && Y == 52) begin oled_data = 16'h64a9; end
    else if (X == 91 && Y == 52) begin oled_data = 16'h64a9; end
    else if (X == 92 && Y == 52) begin oled_data = 16'h64a9; end
    else if (X == 93 && Y == 52) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 52) begin oled_data = 16'h64a9; end
    else if (X == 95 && Y == 52) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 53) begin oled_data = 16'hce16; end
    else if (X == 1 && Y == 53) begin oled_data = 16'h848c; end
    else if (X == 2 && Y == 53) begin oled_data = 16'h53c7; end
    else if (X == 3 && Y == 53) begin oled_data = 16'h6468; end
    else if (X == 4 && Y == 53) begin oled_data = 16'h64a9; end
    else if (X == 5 && Y == 53) begin oled_data = 16'h6468; end
    else if (X == 6 && Y == 53) begin oled_data = 16'h6468; end
    else if (X >= 7 && X <= 8 && Y == 53) begin oled_data = 16'h5c27; end
    else if (X == 9 && Y == 53) begin oled_data = 16'h6468; end
    else if (X == 10 && Y == 53) begin oled_data = 16'h53c7; end
    else if (X == 11 && Y == 53) begin oled_data = 16'hcdd1; end
    else if (X == 13 && Y == 53) begin oled_data = 16'hb550; end
    else if (X == 15 && Y == 53) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 53) begin oled_data = 16'h840f; end
    else if (X >= 17 && X <= 37 && Y == 53) begin oled_data = 16'hcdd1; end
    else if (X == 42 && Y == 53) begin oled_data = 16'hde75; end
    else if (X == 47 && Y == 53) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 53) begin oled_data = 16'had31; end
    else if (X == 57 && Y == 53) begin oled_data = 16'hde75; end
    else if (X >= 61 && X <= 65 && Y == 53) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 53) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 53) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 53) begin oled_data = 16'hb550; end
    else if (X >= 85 && X <= 87 && Y == 53) begin oled_data = 16'hcdd1; end
    else if (X == 88 && Y == 53) begin oled_data = 16'h53c7; end
    else if (X == 89 && Y == 53) begin oled_data = 16'h4346; end
    else if (X == 90 && Y == 53) begin oled_data = 16'h5c27; end
    else if (X == 91 && Y == 53) begin oled_data = 16'h64a9; end
    else if (X == 92 && Y == 53) begin oled_data = 16'h6468; end
    else if (X == 93 && Y == 53) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 53) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 53) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 54) begin oled_data = 16'hce16; end
    else if (X == 3 && Y == 54) begin oled_data = 16'hc5d3; end
    else if (X == 4 && Y == 54) begin oled_data = 16'hb550; end
    else if (X == 5 && Y == 54) begin oled_data = 16'had31; end
    else if (X == 6 && Y == 54) begin oled_data = 16'hb550; end
    else if (X == 7 && Y == 54) begin oled_data = 16'had0f; end
    else if (X == 8 && Y == 54) begin oled_data = 16'ha4ee; end
    else if (X == 9 && Y == 54) begin oled_data = 16'h848c; end
    else if (X == 10 && Y == 54) begin oled_data = 16'h740a; end
    else if (X == 11 && Y == 54) begin oled_data = 16'hb550; end
    else if (X == 13 && Y == 54) begin oled_data = 16'hb550; end
    else if (X >= 14 && X <= 15 && Y == 54) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 54) begin oled_data = 16'h8c71; end
    else if (X >= 18 && X <= 23 && Y == 54) begin oled_data = 16'hcdd1; end
    else if (X == 29 && Y == 54) begin oled_data = 16'hbd91; end
    else if (X >= 30 && X <= 37 && Y == 54) begin oled_data = 16'hcdd1; end
    else if (X == 47 && Y == 54) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 54) begin oled_data = 16'had31; end
    else if (X >= 50 && X <= 75 && Y == 54) begin oled_data = 16'hcdd1; end
    else if (X == 76 && Y == 54) begin oled_data = 16'hcd8f; end
    else if (X == 77 && Y == 54) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 54) begin oled_data = 16'h840f; end
    else if (X == 82 && Y == 54) begin oled_data = 16'hb550; end
    else if (X == 84 && Y == 54) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 54) begin oled_data = 16'ha4f0; end
    else if (X == 87 && Y == 54) begin oled_data = 16'ha4ee; end
    else if (X == 88 && Y == 54) begin oled_data = 16'h3263; end
    else if (X == 89 && Y == 54) begin oled_data = 16'h3b02; end
    else if (X == 90 && Y == 54) begin oled_data = 16'h3b02; end
    else if (X == 91 && Y == 54) begin oled_data = 16'h5c27; end
    else if (X == 92 && Y == 54) begin oled_data = 16'h6468; end
    else if (X >= 93 && X <= 94 && Y == 54) begin oled_data = 16'h5c27; end
    else if (X == 95 && Y == 54) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 55) begin oled_data = 16'hce16; end
    else if (X == 3 && Y == 55) begin oled_data = 16'hde75; end
    else if (X == 4 && Y == 55) begin oled_data = 16'hde75; end
    else if (X == 9 && Y == 55) begin oled_data = 16'hcdd1; end
    else if (X == 13 && Y == 55) begin oled_data = 16'hb550; end
    else if (X == 15 && Y == 55) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 55) begin oled_data = 16'h8c71; end
    else if (X >= 18 && X <= 42 && Y == 55) begin oled_data = 16'hcdd1; end
    else if (X == 47 && Y == 55) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 55) begin oled_data = 16'had31; end
    else if (X >= 50 && X <= 76 && Y == 55) begin oled_data = 16'hcdd1; end
    else if (X == 77 && Y == 55) begin oled_data = 16'hcd8f; end
    else if (X == 78 && Y == 55) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 55) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 55) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 55) begin oled_data = 16'hb550; end
    else if (X == 85 && Y == 55) begin oled_data = 16'hb550; end
    else if (X == 87 && Y == 55) begin oled_data = 16'h7c4b; end
    else if (X == 88 && Y == 55) begin oled_data = 16'h32c3; end
    else if (X == 89 && Y == 55) begin oled_data = 16'h3b02; end
    else if (X == 90 && Y == 55) begin oled_data = 16'h32c3; end
    else if (X == 91 && Y == 55) begin oled_data = 16'h4346; end
    else if (X >= 92 && X <= 94 && Y == 55) begin oled_data = 16'h5c27; end
    else if (X == 95 && Y == 55) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 56) begin oled_data = 16'hb5b6; end
    else if (X == 1 && Y == 56) begin oled_data = 16'h948d; end
    else if (X == 2 && Y == 56) begin oled_data = 16'h848c; end
    else if (X == 3 && Y == 56) begin oled_data = 16'h848c; end
    else if (X == 4 && Y == 56) begin oled_data = 16'h848c; end
    else if (X == 5 && Y == 56) begin oled_data = 16'h740a; end
    else if (X == 6 && Y == 56) begin oled_data = 16'h948d; end
    else if (X == 7 && Y == 56) begin oled_data = 16'had0f; end
    else if (X == 8 && Y == 56) begin oled_data = 16'hbd91; end
    else if (X == 10 && Y == 56) begin oled_data = 16'hcdd1; end
    else if (X == 13 && Y == 56) begin oled_data = 16'had0f; end
    else if (X == 15 && Y == 56) begin oled_data = 16'hbd91; end
    else if (X == 16 && Y == 56) begin oled_data = 16'h8c71; end
    else if (X >= 17 && X <= 24 && Y == 56) begin oled_data = 16'hcdd1; end
    else if (X == 31 && Y == 56) begin oled_data = 16'hbd91; end
    else if (X == 32 && Y == 56) begin oled_data = 16'hbd91; end
    else if (X >= 33 && X <= 43 && Y == 56) begin oled_data = 16'hcdd1; end
    else if (X == 45 && Y == 56) begin oled_data = 16'hbd91; end
    else if (X == 47 && Y == 56) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 56) begin oled_data = 16'ha4f0; end
    else if (X >= 49 && X <= 78 && Y == 56) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 56) begin oled_data = 16'h840f; end
    else if (X == 80 && Y == 56) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 56) begin oled_data = 16'had0f; end
    else if (X == 84 && Y == 56) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 56) begin oled_data = 16'hb550; end
    else if (X == 87 && Y == 56) begin oled_data = 16'had0f; end
    else if (X == 88 && Y == 56) begin oled_data = 16'h2202; end
    else if (X == 89 && Y == 56) begin oled_data = 16'h2202; end
    else if (X == 90 && Y == 56) begin oled_data = 16'h32c3; end
    else if (X == 91 && Y == 56) begin oled_data = 16'h4346; end
    else if (X == 92 && Y == 56) begin oled_data = 16'h53c7; end
    else if (X >= 93 && X <= 94 && Y == 56) begin oled_data = 16'h5c27; end
    else if (X == 95 && Y == 56) begin oled_data = 16'h9551; end
    else if (X == 0 && Y == 57) begin oled_data = 16'hadd4; end
    else if (X == 1 && Y == 57) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 57) begin oled_data = 16'h53c7; end
    else if (X == 3 && Y == 57) begin oled_data = 16'h3263; end
    else if (X == 4 && Y == 57) begin oled_data = 16'h3b02; end
    else if (X == 5 && Y == 57) begin oled_data = 16'h3b02; end
    else if (X == 6 && Y == 57) begin oled_data = 16'h3263; end
    else if (X == 7 && Y == 57) begin oled_data = 16'h4346; end
    else if (X == 8 && Y == 57) begin oled_data = 16'hcdd1; end
    else if (X == 13 && Y == 57) begin oled_data = 16'had0f; end
    else if (X == 15 && Y == 57) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 57) begin oled_data = 16'h840f; end
    else if (X >= 20 && X <= 45 && Y == 57) begin oled_data = 16'hcdd1; end
    else if (X == 47 && Y == 57) begin oled_data = 16'had31; end
    else if (X == 48 && Y == 57) begin oled_data = 16'had31; end
    else if (X >= 49 && X <= 69 && Y == 57) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 57) begin oled_data = 16'h8c71; end
    else if (X == 80 && Y == 57) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 57) begin oled_data = 16'hb550; end
    else if (X == 85 && Y == 57) begin oled_data = 16'hbd91; end
    else if (X == 88 && Y == 57) begin oled_data = 16'h740a; end
    else if (X == 89 && Y == 57) begin oled_data = 16'h53c7; end
    else if (X == 90 && Y == 57) begin oled_data = 16'h5c27; end
    else if (X == 91 && Y == 57) begin oled_data = 16'h6468; end
    else if (X == 92 && Y == 57) begin oled_data = 16'h6468; end
    else if (X == 93 && Y == 57) begin oled_data = 16'h6468; end
    else if (X == 94 && Y == 57) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 57) begin oled_data = 16'h9551; end
    else if (X == 0 && Y == 58) begin oled_data = 16'hadd4; end
    else if (X == 1 && Y == 58) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 58) begin oled_data = 16'h4346; end
    else if (X == 3 && Y == 58) begin oled_data = 16'h2202; end
    else if (X == 4 && Y == 58) begin oled_data = 16'h32c3; end
    else if (X == 5 && Y == 58) begin oled_data = 16'h3263; end
    else if (X == 6 && Y == 58) begin oled_data = 16'h3b02; end
    else if (X == 7 && Y == 58) begin oled_data = 16'h3b02; end
    else if (X == 8 && Y == 58) begin oled_data = 16'h848c; end
    else if (X == 9 && Y == 58) begin oled_data = 16'hcdd1; end
    else if (X == 13 && Y == 58) begin oled_data = 16'had0f; end
    else if (X == 15 && Y == 58) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 58) begin oled_data = 16'h73af; end
    else if (X == 17 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 18 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 19 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 20 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 21 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 22 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 23 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 24 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 25 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 26 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 27 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 28 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 29 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 30 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 31 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 32 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 33 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 34 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 35 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 36 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 37 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 38 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 39 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 40 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 41 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 42 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 43 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 44 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 45 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 46 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 47 && Y == 58) begin oled_data = 16'h840f; end
    else if (X == 48 && Y == 58) begin oled_data = 16'h840f; end
    else if (X == 49 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 50 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 51 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 52 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 53 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 54 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 55 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 56 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 57 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 58 && Y == 58) begin oled_data = 16'h8c71; end
    else if (X == 59 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 60 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 61 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 62 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 63 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 64 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 65 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 66 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 67 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 68 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 69 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 70 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 71 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 72 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 73 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 74 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 75 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 76 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 77 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 78 && Y == 58) begin oled_data = 16'h9cb1; end
    else if (X == 79 && Y == 58) begin oled_data = 16'h73af; end
    else if (X == 80 && Y == 58) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 58) begin oled_data = 16'ha4f0; end
    else if (X == 85 && Y == 58) begin oled_data = 16'hb550; end
    else if (X == 88 && Y == 58) begin oled_data = 16'h63e9; end
    else if (X == 89 && Y == 58) begin oled_data = 16'h5c27; end
    else if (X == 90 && Y == 58) begin oled_data = 16'h6468; end
    else if (X == 91 && Y == 58) begin oled_data = 16'h6468; end
    else if (X == 92 && Y == 58) begin oled_data = 16'h6468; end
    else if (X == 93 && Y == 58) begin oled_data = 16'h5b0c; end
    else if (X == 94 && Y == 58) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 58) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 59) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 59) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 59) begin oled_data = 16'h4346; end
    else if (X == 3 && Y == 59) begin oled_data = 16'h2202; end
    else if (X == 4 && Y == 59) begin oled_data = 16'h3b02; end
    else if (X == 5 && Y == 59) begin oled_data = 16'h3263; end
    else if (X == 6 && Y == 59) begin oled_data = 16'h3263; end
    else if (X == 7 && Y == 59) begin oled_data = 16'h32c3; end
    else if (X == 8 && Y == 59) begin oled_data = 16'h53c7; end
    else if (X == 9 && Y == 59) begin oled_data = 16'h7c4b; end
    else if (X == 10 && Y == 59) begin oled_data = 16'ha4ee; end
    else if (X == 13 && Y == 59) begin oled_data = 16'ha4f0; end
    else if (X == 15 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 16 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 17 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 18 && Y == 59) begin oled_data = 16'hb550; end
    else if (X >= 19 && X <= 20 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 21 && Y == 59) begin oled_data = 16'hb550; end
    else if (X == 22 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 23 && Y == 59) begin oled_data = 16'hb550; end
    else if (X == 24 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 25 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 26 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X >= 27 && X <= 28 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 29 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 30 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 31 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 32 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 33 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 34 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 35 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 36 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 37 && Y == 59) begin oled_data = 16'hb550; end
    else if (X == 38 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 39 && Y == 59) begin oled_data = 16'hb550; end
    else if (X == 40 && Y == 59) begin oled_data = 16'hb550; end
    else if (X == 41 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 42 && Y == 59) begin oled_data = 16'hb550; end
    else if (X == 43 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 44 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 45 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X >= 46 && X <= 49 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 50 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X >= 51 && X <= 52 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 53 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X >= 54 && X <= 55 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 56 && Y == 59) begin oled_data = 16'hc5b2; end
    else if (X == 57 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 58 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X >= 59 && X <= 63 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 64 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 65 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 66 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X >= 67 && X <= 68 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 69 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 70 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 71 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 72 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X >= 73 && X <= 75 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 76 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 77 && Y == 59) begin oled_data = 16'hb550; end
    else if (X == 78 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X == 79 && Y == 59) begin oled_data = 16'hbd91; end
    else if (X >= 80 && X <= 81 && Y == 59) begin oled_data = 16'hcdd1; end
    else if (X == 82 && Y == 59) begin oled_data = 16'had0f; end
    else if (X == 85 && Y == 59) begin oled_data = 16'ha4f0; end
    else if (X == 86 && Y == 59) begin oled_data = 16'h948d; end
    else if (X == 87 && Y == 59) begin oled_data = 16'h740a; end
    else if (X == 88 && Y == 59) begin oled_data = 16'h53c7; end
    else if (X >= 89 && X <= 90 && Y == 59) begin oled_data = 16'h5c27; end
    else if (X == 91 && Y == 59) begin oled_data = 16'h6468; end
    else if (X == 92 && Y == 59) begin oled_data = 16'h4a89; end
    else if (X == 93 && Y == 59) begin oled_data = 16'h622d; end
    else if (X == 94 && Y == 59) begin oled_data = 16'h72ce; end
    else if (X == 95 && Y == 59) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 60) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 60) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 60) begin oled_data = 16'h32c3; end
    else if (X == 3 && Y == 60) begin oled_data = 16'h2202; end
    else if (X == 4 && Y == 60) begin oled_data = 16'h3b02; end
    else if (X == 5 && Y == 60) begin oled_data = 16'h3263; end
    else if (X == 6 && Y == 60) begin oled_data = 16'h2202; end
    else if (X == 7 && Y == 60) begin oled_data = 16'h3263; end
    else if (X >= 8 && X <= 10 && Y == 60) begin oled_data = 16'h5c27; end
    else if (X == 11 && Y == 60) begin oled_data = 16'h740a; end
    else if (X == 12 && Y == 60) begin oled_data = 16'hb550; end
    else if (X == 13 && Y == 60) begin oled_data = 16'h9c8e; end
    else if (X == 18 && Y == 60) begin oled_data = 16'hb550; end
    else if (X >= 23 && X <= 80 && Y == 60) begin oled_data = 16'hcdd1; end
    else if (X == 85 && Y == 60) begin oled_data = 16'h5b88; end
    else if (X == 86 && Y == 60) begin oled_data = 16'h5b0c; end
    else if (X == 87 && Y == 60) begin oled_data = 16'h72ce; end
    else if (X == 88 && Y == 60) begin oled_data = 16'h622d; end
    else if (X == 89 && Y == 60) begin oled_data = 16'h72ce; end
    else if (X == 90 && Y == 60) begin oled_data = 16'h72ce; end
    else if (X == 91 && Y == 60) begin oled_data = 16'h72ce; end
    else if (X == 92 && Y == 60) begin oled_data = 16'h72ce; end
    else if (X == 93 && Y == 60) begin oled_data = 16'h3949; end
    else if (X == 94 && Y == 60) begin oled_data = 16'h3949; end
    else if (X == 95 && Y == 60) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 61) begin oled_data = 16'ha593; end
    else if (X == 1 && Y == 61) begin oled_data = 16'h5c27; end
    else if (X == 2 && Y == 61) begin oled_data = 16'h53c7; end
    else if (X == 3 && Y == 61) begin oled_data = 16'h3263; end
    else if (X == 4 && Y == 61) begin oled_data = 16'h2202; end
    else if (X == 5 && Y == 61) begin oled_data = 16'h32c3; end
    else if (X == 6 && Y == 61) begin oled_data = 16'h4346; end
    else if (X == 7 && Y == 61) begin oled_data = 16'h4346; end
    else if (X >= 8 && X <= 11 && Y == 61) begin oled_data = 16'h5c27; end
    else if (X == 12 && Y == 61) begin oled_data = 16'h53c7; end
    else if (X == 13 && Y == 61) begin oled_data = 16'h4b07; end
    else if (X == 14 && Y == 61) begin oled_data = 16'h5b88; end
    else if (X == 15 && Y == 61) begin oled_data = 16'h5b88; end
    else if (X == 16 && Y == 61) begin oled_data = 16'h5b88; end
    else if (X == 17 && Y == 61) begin oled_data = 16'h5bc8; end
    else if (X == 18 && Y == 61) begin oled_data = 16'h4346; end
    else if (X == 19 && Y == 61) begin oled_data = 16'h5b88; end
    else if (X == 20 && Y == 61) begin oled_data = 16'h948d; end
    else if (X == 21 && Y == 61) begin oled_data = 16'had0f; end
    else if (X == 22 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 23 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 24 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 25 && Y == 61) begin oled_data = 16'hbd91; end
    else if (X == 26 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 27 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 28 && Y == 61) begin oled_data = 16'hbd91; end
    else if (X == 29 && Y == 61) begin oled_data = 16'ha4f0; end
    else if (X == 30 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 31 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 32 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 33 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 34 && Y == 61) begin oled_data = 16'had0f; end
    else if (X == 35 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 36 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 37 && Y == 61) begin oled_data = 16'had0f; end
    else if (X == 38 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 39 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 40 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 41 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 42 && Y == 61) begin oled_data = 16'had0f; end
    else if (X == 43 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 44 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 45 && Y == 61) begin oled_data = 16'had0f; end
    else if (X == 46 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 47 && Y == 61) begin oled_data = 16'ha4f0; end
    else if (X == 48 && Y == 61) begin oled_data = 16'ha4f0; end
    else if (X == 49 && Y == 61) begin oled_data = 16'hbd91; end
    else if (X == 50 && Y == 61) begin oled_data = 16'had0f; end
    else if (X == 51 && Y == 61) begin oled_data = 16'hbd91; end
    else if (X == 52 && Y == 61) begin oled_data = 16'hbd91; end
    else if (X == 53 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 54 && Y == 61) begin oled_data = 16'hbd91; end
    else if (X == 55 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 56 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 57 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 58 && Y == 61) begin oled_data = 16'had0f; end
    else if (X >= 59 && X <= 68 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 69 && Y == 61) begin oled_data = 16'had0f; end
    else if (X == 70 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 71 && Y == 61) begin oled_data = 16'had0f; end
    else if (X == 72 && Y == 61) begin oled_data = 16'had0f; end
    else if (X == 73 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 74 && Y == 61) begin oled_data = 16'had0f; end
    else if (X == 75 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 76 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 77 && Y == 61) begin oled_data = 16'had0f; end
    else if (X == 78 && Y == 61) begin oled_data = 16'had0f; end
    else if (X == 79 && Y == 61) begin oled_data = 16'hb550; end
    else if (X == 80 && Y == 61) begin oled_data = 16'h940c; end
    else if (X == 81 && Y == 61) begin oled_data = 16'h72ce; end
    else if (X == 82 && Y == 61) begin oled_data = 16'h622d; end
    else if (X == 83 && Y == 61) begin oled_data = 16'h72ce; end
    else if (X == 84 && Y == 61) begin oled_data = 16'h622d; end
    else if (X == 85 && Y == 61) begin oled_data = 16'h622d; end
    else if (X == 86 && Y == 61) begin oled_data = 16'h622d; end
    else if (X == 87 && Y == 61) begin oled_data = 16'h622d; end
    else if (X == 88 && Y == 61) begin oled_data = 16'h622d; end
    else if (X == 89 && Y == 61) begin oled_data = 16'h5b0c; end
    else if (X == 90 && Y == 61) begin oled_data = 16'h72ce; end
    else if (X == 91 && Y == 61) begin oled_data = 16'h72ce; end
    else if (X == 92 && Y == 61) begin oled_data = 16'h72ce; end
    else if (X == 93 && Y == 61) begin oled_data = 16'h3949; end
    else if (X == 94 && Y == 61) begin oled_data = 16'h4a89; end
    else if (X == 95 && Y == 61) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 62) begin oled_data = 16'ha593; end
    else if (X >= 1 && X <= 8 && Y == 62) begin oled_data = 16'h5c27; end
    else if (X == 9 && Y == 62) begin oled_data = 16'h6468; end
    else if (X == 10 && Y == 62) begin oled_data = 16'h6468; end
    else if (X == 11 && Y == 62) begin oled_data = 16'h6468; end
    else if (X == 12 && Y == 62) begin oled_data = 16'h6468; end
    else if (X >= 13 && X <= 16 && Y == 62) begin oled_data = 16'h5c27; end
    else if (X == 17 && Y == 62) begin oled_data = 16'h6468; end
    else if (X == 18 && Y == 62) begin oled_data = 16'h6468; end
    else if (X >= 19 && X <= 20 && Y == 62) begin oled_data = 16'h5c27; end
    else if (X == 21 && Y == 62) begin oled_data = 16'h63e9; end
    else if (X == 22 && Y == 62) begin oled_data = 16'h848c; end
    else if (X == 23 && Y == 62) begin oled_data = 16'hb550; end
    else if (X >= 26 && X <= 45 && Y == 62) begin oled_data = 16'hcdd1; end
    else if (X == 46 && Y == 62) begin oled_data = 16'hbd91; end
    else if (X == 47 && Y == 62) begin oled_data = 16'had0f; end
    else if (X == 48 && Y == 62) begin oled_data = 16'hb550; end
    else if (X >= 61 && X <= 77 && Y == 62) begin oled_data = 16'hcdd1; end
    else if (X == 79 && Y == 62) begin oled_data = 16'h9cad; end
    else if (X == 80 && Y == 62) begin oled_data = 16'h53c7; end
    else if (X >= 81 && X <= 83 && Y == 62) begin oled_data = 16'h5c27; end
    else if (X == 84 && Y == 62) begin oled_data = 16'h6468; end
    else if (X == 85 && Y == 62) begin oled_data = 16'h5c27; end
    else if (X == 86 && Y == 62) begin oled_data = 16'h6468; end
    else if (X == 87 && Y == 62) begin oled_data = 16'h6468; end
    else if (X == 88 && Y == 62) begin oled_data = 16'h6468; end
    else if (X == 89 && Y == 62) begin oled_data = 16'h6468; end
    else if (X == 90 && Y == 62) begin oled_data = 16'h6468; end
    else if (X == 91 && Y == 62) begin oled_data = 16'h64a9; end
    else if (X == 92 && Y == 62) begin oled_data = 16'h64a9; end
    else if (X == 93 && Y == 62) begin oled_data = 16'h4b07; end
    else if (X == 94 && Y == 62) begin oled_data = 16'h6468; end
    else if (X == 95 && Y == 62) begin oled_data = 16'ha593; end
    else if (X == 0 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 1 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 2 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 3 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 4 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 5 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 6 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 7 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 8 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 9 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 10 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 11 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 12 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 13 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 14 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 15 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 16 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 17 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 18 && Y == 63) begin oled_data = 16'hadd4; end
    else if (X == 19 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 20 && Y == 63) begin oled_data = 16'hadd4; end
    else if (X == 21 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 22 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 23 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 24 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 25 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 26 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 27 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 28 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 29 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 30 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 31 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 32 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 33 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 34 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 35 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 36 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 37 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 38 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 39 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 40 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 41 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 42 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 43 && Y == 63) begin oled_data = 16'hb573; end
    else if (X == 44 && Y == 63) begin oled_data = 16'h9551; end
    else if (X == 45 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 46 && Y == 63) begin oled_data = 16'h9551; end
    else if (X == 47 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 48 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 49 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 50 && Y == 63) begin oled_data = 16'hb5b6; end
    else if (X == 51 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 52 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 53 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 54 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 55 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 56 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 57 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 58 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 59 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 60 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 61 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 62 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 63 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 64 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 65 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 66 && Y == 63) begin oled_data = 16'hc5d4; end
    else if (X == 67 && Y == 63) begin oled_data = 16'hc5d4; end
    else if (X == 68 && Y == 63) begin oled_data = 16'hc5d4; end
    else if (X == 69 && Y == 63) begin oled_data = 16'hc5d4; end
    else if (X == 70 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 71 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 72 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 73 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 74 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 75 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 76 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 77 && Y == 63) begin oled_data = 16'hce16; end
    else if (X == 78 && Y == 63) begin oled_data = 16'hce57; end
    else if (X == 79 && Y == 63) begin oled_data = 16'hb5b6; end
    else if (X == 80 && Y == 63) begin oled_data = 16'hadd4; end
    else if (X == 81 && Y == 63) begin oled_data = 16'hadd4; end
    else if (X == 82 && Y == 63) begin oled_data = 16'hadd4; end
    else if (X == 83 && Y == 63) begin oled_data = 16'hadd4; end
    else if (X >= 84 && X <= 94 && Y == 63) begin oled_data = 16'ha593; end
    else if (X == 95 && Y == 63) begin oled_data = 16'hce57; end
    else begin oled_data = 16'hd633; end
    
    
    
    end
endmodule
